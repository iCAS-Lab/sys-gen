`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: TODO
// Engineer: TODO
//
// Create Date: 2024-09-06 17:06:52.512677
// Target Devices: TODO
// Tool Versions: TODO
// Description: TODO
//
// Additional Comments:
////////////////////////////////////////////////////////////////////////////////
module mux_1024_to_1 #(parameter SELECT_WIDTH=10, DATA_WIDTH=16) 
(
  input [SELECT_WIDTH-1:0] select,
	input signed [DATA_WIDTH-1:0] in_data_0_0,
	input signed [DATA_WIDTH-1:0] in_data_0_1,
	input signed [DATA_WIDTH-1:0] in_data_0_2,
	input signed [DATA_WIDTH-1:0] in_data_0_3,
	input signed [DATA_WIDTH-1:0] in_data_0_4,
	input signed [DATA_WIDTH-1:0] in_data_0_5,
	input signed [DATA_WIDTH-1:0] in_data_0_6,
	input signed [DATA_WIDTH-1:0] in_data_0_7,
	input signed [DATA_WIDTH-1:0] in_data_0_8,
	input signed [DATA_WIDTH-1:0] in_data_0_9,
	input signed [DATA_WIDTH-1:0] in_data_0_10,
	input signed [DATA_WIDTH-1:0] in_data_0_11,
	input signed [DATA_WIDTH-1:0] in_data_0_12,
	input signed [DATA_WIDTH-1:0] in_data_0_13,
	input signed [DATA_WIDTH-1:0] in_data_0_14,
	input signed [DATA_WIDTH-1:0] in_data_0_15,
	input signed [DATA_WIDTH-1:0] in_data_0_16,
	input signed [DATA_WIDTH-1:0] in_data_0_17,
	input signed [DATA_WIDTH-1:0] in_data_0_18,
	input signed [DATA_WIDTH-1:0] in_data_0_19,
	input signed [DATA_WIDTH-1:0] in_data_0_20,
	input signed [DATA_WIDTH-1:0] in_data_0_21,
	input signed [DATA_WIDTH-1:0] in_data_0_22,
	input signed [DATA_WIDTH-1:0] in_data_0_23,
	input signed [DATA_WIDTH-1:0] in_data_0_24,
	input signed [DATA_WIDTH-1:0] in_data_0_25,
	input signed [DATA_WIDTH-1:0] in_data_0_26,
	input signed [DATA_WIDTH-1:0] in_data_0_27,
	input signed [DATA_WIDTH-1:0] in_data_0_28,
	input signed [DATA_WIDTH-1:0] in_data_0_29,
	input signed [DATA_WIDTH-1:0] in_data_0_30,
	input signed [DATA_WIDTH-1:0] in_data_0_31,
	input signed [DATA_WIDTH-1:0] in_data_1_0,
	input signed [DATA_WIDTH-1:0] in_data_1_1,
	input signed [DATA_WIDTH-1:0] in_data_1_2,
	input signed [DATA_WIDTH-1:0] in_data_1_3,
	input signed [DATA_WIDTH-1:0] in_data_1_4,
	input signed [DATA_WIDTH-1:0] in_data_1_5,
	input signed [DATA_WIDTH-1:0] in_data_1_6,
	input signed [DATA_WIDTH-1:0] in_data_1_7,
	input signed [DATA_WIDTH-1:0] in_data_1_8,
	input signed [DATA_WIDTH-1:0] in_data_1_9,
	input signed [DATA_WIDTH-1:0] in_data_1_10,
	input signed [DATA_WIDTH-1:0] in_data_1_11,
	input signed [DATA_WIDTH-1:0] in_data_1_12,
	input signed [DATA_WIDTH-1:0] in_data_1_13,
	input signed [DATA_WIDTH-1:0] in_data_1_14,
	input signed [DATA_WIDTH-1:0] in_data_1_15,
	input signed [DATA_WIDTH-1:0] in_data_1_16,
	input signed [DATA_WIDTH-1:0] in_data_1_17,
	input signed [DATA_WIDTH-1:0] in_data_1_18,
	input signed [DATA_WIDTH-1:0] in_data_1_19,
	input signed [DATA_WIDTH-1:0] in_data_1_20,
	input signed [DATA_WIDTH-1:0] in_data_1_21,
	input signed [DATA_WIDTH-1:0] in_data_1_22,
	input signed [DATA_WIDTH-1:0] in_data_1_23,
	input signed [DATA_WIDTH-1:0] in_data_1_24,
	input signed [DATA_WIDTH-1:0] in_data_1_25,
	input signed [DATA_WIDTH-1:0] in_data_1_26,
	input signed [DATA_WIDTH-1:0] in_data_1_27,
	input signed [DATA_WIDTH-1:0] in_data_1_28,
	input signed [DATA_WIDTH-1:0] in_data_1_29,
	input signed [DATA_WIDTH-1:0] in_data_1_30,
	input signed [DATA_WIDTH-1:0] in_data_1_31,
	input signed [DATA_WIDTH-1:0] in_data_2_0,
	input signed [DATA_WIDTH-1:0] in_data_2_1,
	input signed [DATA_WIDTH-1:0] in_data_2_2,
	input signed [DATA_WIDTH-1:0] in_data_2_3,
	input signed [DATA_WIDTH-1:0] in_data_2_4,
	input signed [DATA_WIDTH-1:0] in_data_2_5,
	input signed [DATA_WIDTH-1:0] in_data_2_6,
	input signed [DATA_WIDTH-1:0] in_data_2_7,
	input signed [DATA_WIDTH-1:0] in_data_2_8,
	input signed [DATA_WIDTH-1:0] in_data_2_9,
	input signed [DATA_WIDTH-1:0] in_data_2_10,
	input signed [DATA_WIDTH-1:0] in_data_2_11,
	input signed [DATA_WIDTH-1:0] in_data_2_12,
	input signed [DATA_WIDTH-1:0] in_data_2_13,
	input signed [DATA_WIDTH-1:0] in_data_2_14,
	input signed [DATA_WIDTH-1:0] in_data_2_15,
	input signed [DATA_WIDTH-1:0] in_data_2_16,
	input signed [DATA_WIDTH-1:0] in_data_2_17,
	input signed [DATA_WIDTH-1:0] in_data_2_18,
	input signed [DATA_WIDTH-1:0] in_data_2_19,
	input signed [DATA_WIDTH-1:0] in_data_2_20,
	input signed [DATA_WIDTH-1:0] in_data_2_21,
	input signed [DATA_WIDTH-1:0] in_data_2_22,
	input signed [DATA_WIDTH-1:0] in_data_2_23,
	input signed [DATA_WIDTH-1:0] in_data_2_24,
	input signed [DATA_WIDTH-1:0] in_data_2_25,
	input signed [DATA_WIDTH-1:0] in_data_2_26,
	input signed [DATA_WIDTH-1:0] in_data_2_27,
	input signed [DATA_WIDTH-1:0] in_data_2_28,
	input signed [DATA_WIDTH-1:0] in_data_2_29,
	input signed [DATA_WIDTH-1:0] in_data_2_30,
	input signed [DATA_WIDTH-1:0] in_data_2_31,
	input signed [DATA_WIDTH-1:0] in_data_3_0,
	input signed [DATA_WIDTH-1:0] in_data_3_1,
	input signed [DATA_WIDTH-1:0] in_data_3_2,
	input signed [DATA_WIDTH-1:0] in_data_3_3,
	input signed [DATA_WIDTH-1:0] in_data_3_4,
	input signed [DATA_WIDTH-1:0] in_data_3_5,
	input signed [DATA_WIDTH-1:0] in_data_3_6,
	input signed [DATA_WIDTH-1:0] in_data_3_7,
	input signed [DATA_WIDTH-1:0] in_data_3_8,
	input signed [DATA_WIDTH-1:0] in_data_3_9,
	input signed [DATA_WIDTH-1:0] in_data_3_10,
	input signed [DATA_WIDTH-1:0] in_data_3_11,
	input signed [DATA_WIDTH-1:0] in_data_3_12,
	input signed [DATA_WIDTH-1:0] in_data_3_13,
	input signed [DATA_WIDTH-1:0] in_data_3_14,
	input signed [DATA_WIDTH-1:0] in_data_3_15,
	input signed [DATA_WIDTH-1:0] in_data_3_16,
	input signed [DATA_WIDTH-1:0] in_data_3_17,
	input signed [DATA_WIDTH-1:0] in_data_3_18,
	input signed [DATA_WIDTH-1:0] in_data_3_19,
	input signed [DATA_WIDTH-1:0] in_data_3_20,
	input signed [DATA_WIDTH-1:0] in_data_3_21,
	input signed [DATA_WIDTH-1:0] in_data_3_22,
	input signed [DATA_WIDTH-1:0] in_data_3_23,
	input signed [DATA_WIDTH-1:0] in_data_3_24,
	input signed [DATA_WIDTH-1:0] in_data_3_25,
	input signed [DATA_WIDTH-1:0] in_data_3_26,
	input signed [DATA_WIDTH-1:0] in_data_3_27,
	input signed [DATA_WIDTH-1:0] in_data_3_28,
	input signed [DATA_WIDTH-1:0] in_data_3_29,
	input signed [DATA_WIDTH-1:0] in_data_3_30,
	input signed [DATA_WIDTH-1:0] in_data_3_31,
	input signed [DATA_WIDTH-1:0] in_data_4_0,
	input signed [DATA_WIDTH-1:0] in_data_4_1,
	input signed [DATA_WIDTH-1:0] in_data_4_2,
	input signed [DATA_WIDTH-1:0] in_data_4_3,
	input signed [DATA_WIDTH-1:0] in_data_4_4,
	input signed [DATA_WIDTH-1:0] in_data_4_5,
	input signed [DATA_WIDTH-1:0] in_data_4_6,
	input signed [DATA_WIDTH-1:0] in_data_4_7,
	input signed [DATA_WIDTH-1:0] in_data_4_8,
	input signed [DATA_WIDTH-1:0] in_data_4_9,
	input signed [DATA_WIDTH-1:0] in_data_4_10,
	input signed [DATA_WIDTH-1:0] in_data_4_11,
	input signed [DATA_WIDTH-1:0] in_data_4_12,
	input signed [DATA_WIDTH-1:0] in_data_4_13,
	input signed [DATA_WIDTH-1:0] in_data_4_14,
	input signed [DATA_WIDTH-1:0] in_data_4_15,
	input signed [DATA_WIDTH-1:0] in_data_4_16,
	input signed [DATA_WIDTH-1:0] in_data_4_17,
	input signed [DATA_WIDTH-1:0] in_data_4_18,
	input signed [DATA_WIDTH-1:0] in_data_4_19,
	input signed [DATA_WIDTH-1:0] in_data_4_20,
	input signed [DATA_WIDTH-1:0] in_data_4_21,
	input signed [DATA_WIDTH-1:0] in_data_4_22,
	input signed [DATA_WIDTH-1:0] in_data_4_23,
	input signed [DATA_WIDTH-1:0] in_data_4_24,
	input signed [DATA_WIDTH-1:0] in_data_4_25,
	input signed [DATA_WIDTH-1:0] in_data_4_26,
	input signed [DATA_WIDTH-1:0] in_data_4_27,
	input signed [DATA_WIDTH-1:0] in_data_4_28,
	input signed [DATA_WIDTH-1:0] in_data_4_29,
	input signed [DATA_WIDTH-1:0] in_data_4_30,
	input signed [DATA_WIDTH-1:0] in_data_4_31,
	input signed [DATA_WIDTH-1:0] in_data_5_0,
	input signed [DATA_WIDTH-1:0] in_data_5_1,
	input signed [DATA_WIDTH-1:0] in_data_5_2,
	input signed [DATA_WIDTH-1:0] in_data_5_3,
	input signed [DATA_WIDTH-1:0] in_data_5_4,
	input signed [DATA_WIDTH-1:0] in_data_5_5,
	input signed [DATA_WIDTH-1:0] in_data_5_6,
	input signed [DATA_WIDTH-1:0] in_data_5_7,
	input signed [DATA_WIDTH-1:0] in_data_5_8,
	input signed [DATA_WIDTH-1:0] in_data_5_9,
	input signed [DATA_WIDTH-1:0] in_data_5_10,
	input signed [DATA_WIDTH-1:0] in_data_5_11,
	input signed [DATA_WIDTH-1:0] in_data_5_12,
	input signed [DATA_WIDTH-1:0] in_data_5_13,
	input signed [DATA_WIDTH-1:0] in_data_5_14,
	input signed [DATA_WIDTH-1:0] in_data_5_15,
	input signed [DATA_WIDTH-1:0] in_data_5_16,
	input signed [DATA_WIDTH-1:0] in_data_5_17,
	input signed [DATA_WIDTH-1:0] in_data_5_18,
	input signed [DATA_WIDTH-1:0] in_data_5_19,
	input signed [DATA_WIDTH-1:0] in_data_5_20,
	input signed [DATA_WIDTH-1:0] in_data_5_21,
	input signed [DATA_WIDTH-1:0] in_data_5_22,
	input signed [DATA_WIDTH-1:0] in_data_5_23,
	input signed [DATA_WIDTH-1:0] in_data_5_24,
	input signed [DATA_WIDTH-1:0] in_data_5_25,
	input signed [DATA_WIDTH-1:0] in_data_5_26,
	input signed [DATA_WIDTH-1:0] in_data_5_27,
	input signed [DATA_WIDTH-1:0] in_data_5_28,
	input signed [DATA_WIDTH-1:0] in_data_5_29,
	input signed [DATA_WIDTH-1:0] in_data_5_30,
	input signed [DATA_WIDTH-1:0] in_data_5_31,
	input signed [DATA_WIDTH-1:0] in_data_6_0,
	input signed [DATA_WIDTH-1:0] in_data_6_1,
	input signed [DATA_WIDTH-1:0] in_data_6_2,
	input signed [DATA_WIDTH-1:0] in_data_6_3,
	input signed [DATA_WIDTH-1:0] in_data_6_4,
	input signed [DATA_WIDTH-1:0] in_data_6_5,
	input signed [DATA_WIDTH-1:0] in_data_6_6,
	input signed [DATA_WIDTH-1:0] in_data_6_7,
	input signed [DATA_WIDTH-1:0] in_data_6_8,
	input signed [DATA_WIDTH-1:0] in_data_6_9,
	input signed [DATA_WIDTH-1:0] in_data_6_10,
	input signed [DATA_WIDTH-1:0] in_data_6_11,
	input signed [DATA_WIDTH-1:0] in_data_6_12,
	input signed [DATA_WIDTH-1:0] in_data_6_13,
	input signed [DATA_WIDTH-1:0] in_data_6_14,
	input signed [DATA_WIDTH-1:0] in_data_6_15,
	input signed [DATA_WIDTH-1:0] in_data_6_16,
	input signed [DATA_WIDTH-1:0] in_data_6_17,
	input signed [DATA_WIDTH-1:0] in_data_6_18,
	input signed [DATA_WIDTH-1:0] in_data_6_19,
	input signed [DATA_WIDTH-1:0] in_data_6_20,
	input signed [DATA_WIDTH-1:0] in_data_6_21,
	input signed [DATA_WIDTH-1:0] in_data_6_22,
	input signed [DATA_WIDTH-1:0] in_data_6_23,
	input signed [DATA_WIDTH-1:0] in_data_6_24,
	input signed [DATA_WIDTH-1:0] in_data_6_25,
	input signed [DATA_WIDTH-1:0] in_data_6_26,
	input signed [DATA_WIDTH-1:0] in_data_6_27,
	input signed [DATA_WIDTH-1:0] in_data_6_28,
	input signed [DATA_WIDTH-1:0] in_data_6_29,
	input signed [DATA_WIDTH-1:0] in_data_6_30,
	input signed [DATA_WIDTH-1:0] in_data_6_31,
	input signed [DATA_WIDTH-1:0] in_data_7_0,
	input signed [DATA_WIDTH-1:0] in_data_7_1,
	input signed [DATA_WIDTH-1:0] in_data_7_2,
	input signed [DATA_WIDTH-1:0] in_data_7_3,
	input signed [DATA_WIDTH-1:0] in_data_7_4,
	input signed [DATA_WIDTH-1:0] in_data_7_5,
	input signed [DATA_WIDTH-1:0] in_data_7_6,
	input signed [DATA_WIDTH-1:0] in_data_7_7,
	input signed [DATA_WIDTH-1:0] in_data_7_8,
	input signed [DATA_WIDTH-1:0] in_data_7_9,
	input signed [DATA_WIDTH-1:0] in_data_7_10,
	input signed [DATA_WIDTH-1:0] in_data_7_11,
	input signed [DATA_WIDTH-1:0] in_data_7_12,
	input signed [DATA_WIDTH-1:0] in_data_7_13,
	input signed [DATA_WIDTH-1:0] in_data_7_14,
	input signed [DATA_WIDTH-1:0] in_data_7_15,
	input signed [DATA_WIDTH-1:0] in_data_7_16,
	input signed [DATA_WIDTH-1:0] in_data_7_17,
	input signed [DATA_WIDTH-1:0] in_data_7_18,
	input signed [DATA_WIDTH-1:0] in_data_7_19,
	input signed [DATA_WIDTH-1:0] in_data_7_20,
	input signed [DATA_WIDTH-1:0] in_data_7_21,
	input signed [DATA_WIDTH-1:0] in_data_7_22,
	input signed [DATA_WIDTH-1:0] in_data_7_23,
	input signed [DATA_WIDTH-1:0] in_data_7_24,
	input signed [DATA_WIDTH-1:0] in_data_7_25,
	input signed [DATA_WIDTH-1:0] in_data_7_26,
	input signed [DATA_WIDTH-1:0] in_data_7_27,
	input signed [DATA_WIDTH-1:0] in_data_7_28,
	input signed [DATA_WIDTH-1:0] in_data_7_29,
	input signed [DATA_WIDTH-1:0] in_data_7_30,
	input signed [DATA_WIDTH-1:0] in_data_7_31,
	input signed [DATA_WIDTH-1:0] in_data_8_0,
	input signed [DATA_WIDTH-1:0] in_data_8_1,
	input signed [DATA_WIDTH-1:0] in_data_8_2,
	input signed [DATA_WIDTH-1:0] in_data_8_3,
	input signed [DATA_WIDTH-1:0] in_data_8_4,
	input signed [DATA_WIDTH-1:0] in_data_8_5,
	input signed [DATA_WIDTH-1:0] in_data_8_6,
	input signed [DATA_WIDTH-1:0] in_data_8_7,
	input signed [DATA_WIDTH-1:0] in_data_8_8,
	input signed [DATA_WIDTH-1:0] in_data_8_9,
	input signed [DATA_WIDTH-1:0] in_data_8_10,
	input signed [DATA_WIDTH-1:0] in_data_8_11,
	input signed [DATA_WIDTH-1:0] in_data_8_12,
	input signed [DATA_WIDTH-1:0] in_data_8_13,
	input signed [DATA_WIDTH-1:0] in_data_8_14,
	input signed [DATA_WIDTH-1:0] in_data_8_15,
	input signed [DATA_WIDTH-1:0] in_data_8_16,
	input signed [DATA_WIDTH-1:0] in_data_8_17,
	input signed [DATA_WIDTH-1:0] in_data_8_18,
	input signed [DATA_WIDTH-1:0] in_data_8_19,
	input signed [DATA_WIDTH-1:0] in_data_8_20,
	input signed [DATA_WIDTH-1:0] in_data_8_21,
	input signed [DATA_WIDTH-1:0] in_data_8_22,
	input signed [DATA_WIDTH-1:0] in_data_8_23,
	input signed [DATA_WIDTH-1:0] in_data_8_24,
	input signed [DATA_WIDTH-1:0] in_data_8_25,
	input signed [DATA_WIDTH-1:0] in_data_8_26,
	input signed [DATA_WIDTH-1:0] in_data_8_27,
	input signed [DATA_WIDTH-1:0] in_data_8_28,
	input signed [DATA_WIDTH-1:0] in_data_8_29,
	input signed [DATA_WIDTH-1:0] in_data_8_30,
	input signed [DATA_WIDTH-1:0] in_data_8_31,
	input signed [DATA_WIDTH-1:0] in_data_9_0,
	input signed [DATA_WIDTH-1:0] in_data_9_1,
	input signed [DATA_WIDTH-1:0] in_data_9_2,
	input signed [DATA_WIDTH-1:0] in_data_9_3,
	input signed [DATA_WIDTH-1:0] in_data_9_4,
	input signed [DATA_WIDTH-1:0] in_data_9_5,
	input signed [DATA_WIDTH-1:0] in_data_9_6,
	input signed [DATA_WIDTH-1:0] in_data_9_7,
	input signed [DATA_WIDTH-1:0] in_data_9_8,
	input signed [DATA_WIDTH-1:0] in_data_9_9,
	input signed [DATA_WIDTH-1:0] in_data_9_10,
	input signed [DATA_WIDTH-1:0] in_data_9_11,
	input signed [DATA_WIDTH-1:0] in_data_9_12,
	input signed [DATA_WIDTH-1:0] in_data_9_13,
	input signed [DATA_WIDTH-1:0] in_data_9_14,
	input signed [DATA_WIDTH-1:0] in_data_9_15,
	input signed [DATA_WIDTH-1:0] in_data_9_16,
	input signed [DATA_WIDTH-1:0] in_data_9_17,
	input signed [DATA_WIDTH-1:0] in_data_9_18,
	input signed [DATA_WIDTH-1:0] in_data_9_19,
	input signed [DATA_WIDTH-1:0] in_data_9_20,
	input signed [DATA_WIDTH-1:0] in_data_9_21,
	input signed [DATA_WIDTH-1:0] in_data_9_22,
	input signed [DATA_WIDTH-1:0] in_data_9_23,
	input signed [DATA_WIDTH-1:0] in_data_9_24,
	input signed [DATA_WIDTH-1:0] in_data_9_25,
	input signed [DATA_WIDTH-1:0] in_data_9_26,
	input signed [DATA_WIDTH-1:0] in_data_9_27,
	input signed [DATA_WIDTH-1:0] in_data_9_28,
	input signed [DATA_WIDTH-1:0] in_data_9_29,
	input signed [DATA_WIDTH-1:0] in_data_9_30,
	input signed [DATA_WIDTH-1:0] in_data_9_31,
	input signed [DATA_WIDTH-1:0] in_data_10_0,
	input signed [DATA_WIDTH-1:0] in_data_10_1,
	input signed [DATA_WIDTH-1:0] in_data_10_2,
	input signed [DATA_WIDTH-1:0] in_data_10_3,
	input signed [DATA_WIDTH-1:0] in_data_10_4,
	input signed [DATA_WIDTH-1:0] in_data_10_5,
	input signed [DATA_WIDTH-1:0] in_data_10_6,
	input signed [DATA_WIDTH-1:0] in_data_10_7,
	input signed [DATA_WIDTH-1:0] in_data_10_8,
	input signed [DATA_WIDTH-1:0] in_data_10_9,
	input signed [DATA_WIDTH-1:0] in_data_10_10,
	input signed [DATA_WIDTH-1:0] in_data_10_11,
	input signed [DATA_WIDTH-1:0] in_data_10_12,
	input signed [DATA_WIDTH-1:0] in_data_10_13,
	input signed [DATA_WIDTH-1:0] in_data_10_14,
	input signed [DATA_WIDTH-1:0] in_data_10_15,
	input signed [DATA_WIDTH-1:0] in_data_10_16,
	input signed [DATA_WIDTH-1:0] in_data_10_17,
	input signed [DATA_WIDTH-1:0] in_data_10_18,
	input signed [DATA_WIDTH-1:0] in_data_10_19,
	input signed [DATA_WIDTH-1:0] in_data_10_20,
	input signed [DATA_WIDTH-1:0] in_data_10_21,
	input signed [DATA_WIDTH-1:0] in_data_10_22,
	input signed [DATA_WIDTH-1:0] in_data_10_23,
	input signed [DATA_WIDTH-1:0] in_data_10_24,
	input signed [DATA_WIDTH-1:0] in_data_10_25,
	input signed [DATA_WIDTH-1:0] in_data_10_26,
	input signed [DATA_WIDTH-1:0] in_data_10_27,
	input signed [DATA_WIDTH-1:0] in_data_10_28,
	input signed [DATA_WIDTH-1:0] in_data_10_29,
	input signed [DATA_WIDTH-1:0] in_data_10_30,
	input signed [DATA_WIDTH-1:0] in_data_10_31,
	input signed [DATA_WIDTH-1:0] in_data_11_0,
	input signed [DATA_WIDTH-1:0] in_data_11_1,
	input signed [DATA_WIDTH-1:0] in_data_11_2,
	input signed [DATA_WIDTH-1:0] in_data_11_3,
	input signed [DATA_WIDTH-1:0] in_data_11_4,
	input signed [DATA_WIDTH-1:0] in_data_11_5,
	input signed [DATA_WIDTH-1:0] in_data_11_6,
	input signed [DATA_WIDTH-1:0] in_data_11_7,
	input signed [DATA_WIDTH-1:0] in_data_11_8,
	input signed [DATA_WIDTH-1:0] in_data_11_9,
	input signed [DATA_WIDTH-1:0] in_data_11_10,
	input signed [DATA_WIDTH-1:0] in_data_11_11,
	input signed [DATA_WIDTH-1:0] in_data_11_12,
	input signed [DATA_WIDTH-1:0] in_data_11_13,
	input signed [DATA_WIDTH-1:0] in_data_11_14,
	input signed [DATA_WIDTH-1:0] in_data_11_15,
	input signed [DATA_WIDTH-1:0] in_data_11_16,
	input signed [DATA_WIDTH-1:0] in_data_11_17,
	input signed [DATA_WIDTH-1:0] in_data_11_18,
	input signed [DATA_WIDTH-1:0] in_data_11_19,
	input signed [DATA_WIDTH-1:0] in_data_11_20,
	input signed [DATA_WIDTH-1:0] in_data_11_21,
	input signed [DATA_WIDTH-1:0] in_data_11_22,
	input signed [DATA_WIDTH-1:0] in_data_11_23,
	input signed [DATA_WIDTH-1:0] in_data_11_24,
	input signed [DATA_WIDTH-1:0] in_data_11_25,
	input signed [DATA_WIDTH-1:0] in_data_11_26,
	input signed [DATA_WIDTH-1:0] in_data_11_27,
	input signed [DATA_WIDTH-1:0] in_data_11_28,
	input signed [DATA_WIDTH-1:0] in_data_11_29,
	input signed [DATA_WIDTH-1:0] in_data_11_30,
	input signed [DATA_WIDTH-1:0] in_data_11_31,
	input signed [DATA_WIDTH-1:0] in_data_12_0,
	input signed [DATA_WIDTH-1:0] in_data_12_1,
	input signed [DATA_WIDTH-1:0] in_data_12_2,
	input signed [DATA_WIDTH-1:0] in_data_12_3,
	input signed [DATA_WIDTH-1:0] in_data_12_4,
	input signed [DATA_WIDTH-1:0] in_data_12_5,
	input signed [DATA_WIDTH-1:0] in_data_12_6,
	input signed [DATA_WIDTH-1:0] in_data_12_7,
	input signed [DATA_WIDTH-1:0] in_data_12_8,
	input signed [DATA_WIDTH-1:0] in_data_12_9,
	input signed [DATA_WIDTH-1:0] in_data_12_10,
	input signed [DATA_WIDTH-1:0] in_data_12_11,
	input signed [DATA_WIDTH-1:0] in_data_12_12,
	input signed [DATA_WIDTH-1:0] in_data_12_13,
	input signed [DATA_WIDTH-1:0] in_data_12_14,
	input signed [DATA_WIDTH-1:0] in_data_12_15,
	input signed [DATA_WIDTH-1:0] in_data_12_16,
	input signed [DATA_WIDTH-1:0] in_data_12_17,
	input signed [DATA_WIDTH-1:0] in_data_12_18,
	input signed [DATA_WIDTH-1:0] in_data_12_19,
	input signed [DATA_WIDTH-1:0] in_data_12_20,
	input signed [DATA_WIDTH-1:0] in_data_12_21,
	input signed [DATA_WIDTH-1:0] in_data_12_22,
	input signed [DATA_WIDTH-1:0] in_data_12_23,
	input signed [DATA_WIDTH-1:0] in_data_12_24,
	input signed [DATA_WIDTH-1:0] in_data_12_25,
	input signed [DATA_WIDTH-1:0] in_data_12_26,
	input signed [DATA_WIDTH-1:0] in_data_12_27,
	input signed [DATA_WIDTH-1:0] in_data_12_28,
	input signed [DATA_WIDTH-1:0] in_data_12_29,
	input signed [DATA_WIDTH-1:0] in_data_12_30,
	input signed [DATA_WIDTH-1:0] in_data_12_31,
	input signed [DATA_WIDTH-1:0] in_data_13_0,
	input signed [DATA_WIDTH-1:0] in_data_13_1,
	input signed [DATA_WIDTH-1:0] in_data_13_2,
	input signed [DATA_WIDTH-1:0] in_data_13_3,
	input signed [DATA_WIDTH-1:0] in_data_13_4,
	input signed [DATA_WIDTH-1:0] in_data_13_5,
	input signed [DATA_WIDTH-1:0] in_data_13_6,
	input signed [DATA_WIDTH-1:0] in_data_13_7,
	input signed [DATA_WIDTH-1:0] in_data_13_8,
	input signed [DATA_WIDTH-1:0] in_data_13_9,
	input signed [DATA_WIDTH-1:0] in_data_13_10,
	input signed [DATA_WIDTH-1:0] in_data_13_11,
	input signed [DATA_WIDTH-1:0] in_data_13_12,
	input signed [DATA_WIDTH-1:0] in_data_13_13,
	input signed [DATA_WIDTH-1:0] in_data_13_14,
	input signed [DATA_WIDTH-1:0] in_data_13_15,
	input signed [DATA_WIDTH-1:0] in_data_13_16,
	input signed [DATA_WIDTH-1:0] in_data_13_17,
	input signed [DATA_WIDTH-1:0] in_data_13_18,
	input signed [DATA_WIDTH-1:0] in_data_13_19,
	input signed [DATA_WIDTH-1:0] in_data_13_20,
	input signed [DATA_WIDTH-1:0] in_data_13_21,
	input signed [DATA_WIDTH-1:0] in_data_13_22,
	input signed [DATA_WIDTH-1:0] in_data_13_23,
	input signed [DATA_WIDTH-1:0] in_data_13_24,
	input signed [DATA_WIDTH-1:0] in_data_13_25,
	input signed [DATA_WIDTH-1:0] in_data_13_26,
	input signed [DATA_WIDTH-1:0] in_data_13_27,
	input signed [DATA_WIDTH-1:0] in_data_13_28,
	input signed [DATA_WIDTH-1:0] in_data_13_29,
	input signed [DATA_WIDTH-1:0] in_data_13_30,
	input signed [DATA_WIDTH-1:0] in_data_13_31,
	input signed [DATA_WIDTH-1:0] in_data_14_0,
	input signed [DATA_WIDTH-1:0] in_data_14_1,
	input signed [DATA_WIDTH-1:0] in_data_14_2,
	input signed [DATA_WIDTH-1:0] in_data_14_3,
	input signed [DATA_WIDTH-1:0] in_data_14_4,
	input signed [DATA_WIDTH-1:0] in_data_14_5,
	input signed [DATA_WIDTH-1:0] in_data_14_6,
	input signed [DATA_WIDTH-1:0] in_data_14_7,
	input signed [DATA_WIDTH-1:0] in_data_14_8,
	input signed [DATA_WIDTH-1:0] in_data_14_9,
	input signed [DATA_WIDTH-1:0] in_data_14_10,
	input signed [DATA_WIDTH-1:0] in_data_14_11,
	input signed [DATA_WIDTH-1:0] in_data_14_12,
	input signed [DATA_WIDTH-1:0] in_data_14_13,
	input signed [DATA_WIDTH-1:0] in_data_14_14,
	input signed [DATA_WIDTH-1:0] in_data_14_15,
	input signed [DATA_WIDTH-1:0] in_data_14_16,
	input signed [DATA_WIDTH-1:0] in_data_14_17,
	input signed [DATA_WIDTH-1:0] in_data_14_18,
	input signed [DATA_WIDTH-1:0] in_data_14_19,
	input signed [DATA_WIDTH-1:0] in_data_14_20,
	input signed [DATA_WIDTH-1:0] in_data_14_21,
	input signed [DATA_WIDTH-1:0] in_data_14_22,
	input signed [DATA_WIDTH-1:0] in_data_14_23,
	input signed [DATA_WIDTH-1:0] in_data_14_24,
	input signed [DATA_WIDTH-1:0] in_data_14_25,
	input signed [DATA_WIDTH-1:0] in_data_14_26,
	input signed [DATA_WIDTH-1:0] in_data_14_27,
	input signed [DATA_WIDTH-1:0] in_data_14_28,
	input signed [DATA_WIDTH-1:0] in_data_14_29,
	input signed [DATA_WIDTH-1:0] in_data_14_30,
	input signed [DATA_WIDTH-1:0] in_data_14_31,
	input signed [DATA_WIDTH-1:0] in_data_15_0,
	input signed [DATA_WIDTH-1:0] in_data_15_1,
	input signed [DATA_WIDTH-1:0] in_data_15_2,
	input signed [DATA_WIDTH-1:0] in_data_15_3,
	input signed [DATA_WIDTH-1:0] in_data_15_4,
	input signed [DATA_WIDTH-1:0] in_data_15_5,
	input signed [DATA_WIDTH-1:0] in_data_15_6,
	input signed [DATA_WIDTH-1:0] in_data_15_7,
	input signed [DATA_WIDTH-1:0] in_data_15_8,
	input signed [DATA_WIDTH-1:0] in_data_15_9,
	input signed [DATA_WIDTH-1:0] in_data_15_10,
	input signed [DATA_WIDTH-1:0] in_data_15_11,
	input signed [DATA_WIDTH-1:0] in_data_15_12,
	input signed [DATA_WIDTH-1:0] in_data_15_13,
	input signed [DATA_WIDTH-1:0] in_data_15_14,
	input signed [DATA_WIDTH-1:0] in_data_15_15,
	input signed [DATA_WIDTH-1:0] in_data_15_16,
	input signed [DATA_WIDTH-1:0] in_data_15_17,
	input signed [DATA_WIDTH-1:0] in_data_15_18,
	input signed [DATA_WIDTH-1:0] in_data_15_19,
	input signed [DATA_WIDTH-1:0] in_data_15_20,
	input signed [DATA_WIDTH-1:0] in_data_15_21,
	input signed [DATA_WIDTH-1:0] in_data_15_22,
	input signed [DATA_WIDTH-1:0] in_data_15_23,
	input signed [DATA_WIDTH-1:0] in_data_15_24,
	input signed [DATA_WIDTH-1:0] in_data_15_25,
	input signed [DATA_WIDTH-1:0] in_data_15_26,
	input signed [DATA_WIDTH-1:0] in_data_15_27,
	input signed [DATA_WIDTH-1:0] in_data_15_28,
	input signed [DATA_WIDTH-1:0] in_data_15_29,
	input signed [DATA_WIDTH-1:0] in_data_15_30,
	input signed [DATA_WIDTH-1:0] in_data_15_31,
	input signed [DATA_WIDTH-1:0] in_data_16_0,
	input signed [DATA_WIDTH-1:0] in_data_16_1,
	input signed [DATA_WIDTH-1:0] in_data_16_2,
	input signed [DATA_WIDTH-1:0] in_data_16_3,
	input signed [DATA_WIDTH-1:0] in_data_16_4,
	input signed [DATA_WIDTH-1:0] in_data_16_5,
	input signed [DATA_WIDTH-1:0] in_data_16_6,
	input signed [DATA_WIDTH-1:0] in_data_16_7,
	input signed [DATA_WIDTH-1:0] in_data_16_8,
	input signed [DATA_WIDTH-1:0] in_data_16_9,
	input signed [DATA_WIDTH-1:0] in_data_16_10,
	input signed [DATA_WIDTH-1:0] in_data_16_11,
	input signed [DATA_WIDTH-1:0] in_data_16_12,
	input signed [DATA_WIDTH-1:0] in_data_16_13,
	input signed [DATA_WIDTH-1:0] in_data_16_14,
	input signed [DATA_WIDTH-1:0] in_data_16_15,
	input signed [DATA_WIDTH-1:0] in_data_16_16,
	input signed [DATA_WIDTH-1:0] in_data_16_17,
	input signed [DATA_WIDTH-1:0] in_data_16_18,
	input signed [DATA_WIDTH-1:0] in_data_16_19,
	input signed [DATA_WIDTH-1:0] in_data_16_20,
	input signed [DATA_WIDTH-1:0] in_data_16_21,
	input signed [DATA_WIDTH-1:0] in_data_16_22,
	input signed [DATA_WIDTH-1:0] in_data_16_23,
	input signed [DATA_WIDTH-1:0] in_data_16_24,
	input signed [DATA_WIDTH-1:0] in_data_16_25,
	input signed [DATA_WIDTH-1:0] in_data_16_26,
	input signed [DATA_WIDTH-1:0] in_data_16_27,
	input signed [DATA_WIDTH-1:0] in_data_16_28,
	input signed [DATA_WIDTH-1:0] in_data_16_29,
	input signed [DATA_WIDTH-1:0] in_data_16_30,
	input signed [DATA_WIDTH-1:0] in_data_16_31,
	input signed [DATA_WIDTH-1:0] in_data_17_0,
	input signed [DATA_WIDTH-1:0] in_data_17_1,
	input signed [DATA_WIDTH-1:0] in_data_17_2,
	input signed [DATA_WIDTH-1:0] in_data_17_3,
	input signed [DATA_WIDTH-1:0] in_data_17_4,
	input signed [DATA_WIDTH-1:0] in_data_17_5,
	input signed [DATA_WIDTH-1:0] in_data_17_6,
	input signed [DATA_WIDTH-1:0] in_data_17_7,
	input signed [DATA_WIDTH-1:0] in_data_17_8,
	input signed [DATA_WIDTH-1:0] in_data_17_9,
	input signed [DATA_WIDTH-1:0] in_data_17_10,
	input signed [DATA_WIDTH-1:0] in_data_17_11,
	input signed [DATA_WIDTH-1:0] in_data_17_12,
	input signed [DATA_WIDTH-1:0] in_data_17_13,
	input signed [DATA_WIDTH-1:0] in_data_17_14,
	input signed [DATA_WIDTH-1:0] in_data_17_15,
	input signed [DATA_WIDTH-1:0] in_data_17_16,
	input signed [DATA_WIDTH-1:0] in_data_17_17,
	input signed [DATA_WIDTH-1:0] in_data_17_18,
	input signed [DATA_WIDTH-1:0] in_data_17_19,
	input signed [DATA_WIDTH-1:0] in_data_17_20,
	input signed [DATA_WIDTH-1:0] in_data_17_21,
	input signed [DATA_WIDTH-1:0] in_data_17_22,
	input signed [DATA_WIDTH-1:0] in_data_17_23,
	input signed [DATA_WIDTH-1:0] in_data_17_24,
	input signed [DATA_WIDTH-1:0] in_data_17_25,
	input signed [DATA_WIDTH-1:0] in_data_17_26,
	input signed [DATA_WIDTH-1:0] in_data_17_27,
	input signed [DATA_WIDTH-1:0] in_data_17_28,
	input signed [DATA_WIDTH-1:0] in_data_17_29,
	input signed [DATA_WIDTH-1:0] in_data_17_30,
	input signed [DATA_WIDTH-1:0] in_data_17_31,
	input signed [DATA_WIDTH-1:0] in_data_18_0,
	input signed [DATA_WIDTH-1:0] in_data_18_1,
	input signed [DATA_WIDTH-1:0] in_data_18_2,
	input signed [DATA_WIDTH-1:0] in_data_18_3,
	input signed [DATA_WIDTH-1:0] in_data_18_4,
	input signed [DATA_WIDTH-1:0] in_data_18_5,
	input signed [DATA_WIDTH-1:0] in_data_18_6,
	input signed [DATA_WIDTH-1:0] in_data_18_7,
	input signed [DATA_WIDTH-1:0] in_data_18_8,
	input signed [DATA_WIDTH-1:0] in_data_18_9,
	input signed [DATA_WIDTH-1:0] in_data_18_10,
	input signed [DATA_WIDTH-1:0] in_data_18_11,
	input signed [DATA_WIDTH-1:0] in_data_18_12,
	input signed [DATA_WIDTH-1:0] in_data_18_13,
	input signed [DATA_WIDTH-1:0] in_data_18_14,
	input signed [DATA_WIDTH-1:0] in_data_18_15,
	input signed [DATA_WIDTH-1:0] in_data_18_16,
	input signed [DATA_WIDTH-1:0] in_data_18_17,
	input signed [DATA_WIDTH-1:0] in_data_18_18,
	input signed [DATA_WIDTH-1:0] in_data_18_19,
	input signed [DATA_WIDTH-1:0] in_data_18_20,
	input signed [DATA_WIDTH-1:0] in_data_18_21,
	input signed [DATA_WIDTH-1:0] in_data_18_22,
	input signed [DATA_WIDTH-1:0] in_data_18_23,
	input signed [DATA_WIDTH-1:0] in_data_18_24,
	input signed [DATA_WIDTH-1:0] in_data_18_25,
	input signed [DATA_WIDTH-1:0] in_data_18_26,
	input signed [DATA_WIDTH-1:0] in_data_18_27,
	input signed [DATA_WIDTH-1:0] in_data_18_28,
	input signed [DATA_WIDTH-1:0] in_data_18_29,
	input signed [DATA_WIDTH-1:0] in_data_18_30,
	input signed [DATA_WIDTH-1:0] in_data_18_31,
	input signed [DATA_WIDTH-1:0] in_data_19_0,
	input signed [DATA_WIDTH-1:0] in_data_19_1,
	input signed [DATA_WIDTH-1:0] in_data_19_2,
	input signed [DATA_WIDTH-1:0] in_data_19_3,
	input signed [DATA_WIDTH-1:0] in_data_19_4,
	input signed [DATA_WIDTH-1:0] in_data_19_5,
	input signed [DATA_WIDTH-1:0] in_data_19_6,
	input signed [DATA_WIDTH-1:0] in_data_19_7,
	input signed [DATA_WIDTH-1:0] in_data_19_8,
	input signed [DATA_WIDTH-1:0] in_data_19_9,
	input signed [DATA_WIDTH-1:0] in_data_19_10,
	input signed [DATA_WIDTH-1:0] in_data_19_11,
	input signed [DATA_WIDTH-1:0] in_data_19_12,
	input signed [DATA_WIDTH-1:0] in_data_19_13,
	input signed [DATA_WIDTH-1:0] in_data_19_14,
	input signed [DATA_WIDTH-1:0] in_data_19_15,
	input signed [DATA_WIDTH-1:0] in_data_19_16,
	input signed [DATA_WIDTH-1:0] in_data_19_17,
	input signed [DATA_WIDTH-1:0] in_data_19_18,
	input signed [DATA_WIDTH-1:0] in_data_19_19,
	input signed [DATA_WIDTH-1:0] in_data_19_20,
	input signed [DATA_WIDTH-1:0] in_data_19_21,
	input signed [DATA_WIDTH-1:0] in_data_19_22,
	input signed [DATA_WIDTH-1:0] in_data_19_23,
	input signed [DATA_WIDTH-1:0] in_data_19_24,
	input signed [DATA_WIDTH-1:0] in_data_19_25,
	input signed [DATA_WIDTH-1:0] in_data_19_26,
	input signed [DATA_WIDTH-1:0] in_data_19_27,
	input signed [DATA_WIDTH-1:0] in_data_19_28,
	input signed [DATA_WIDTH-1:0] in_data_19_29,
	input signed [DATA_WIDTH-1:0] in_data_19_30,
	input signed [DATA_WIDTH-1:0] in_data_19_31,
	input signed [DATA_WIDTH-1:0] in_data_20_0,
	input signed [DATA_WIDTH-1:0] in_data_20_1,
	input signed [DATA_WIDTH-1:0] in_data_20_2,
	input signed [DATA_WIDTH-1:0] in_data_20_3,
	input signed [DATA_WIDTH-1:0] in_data_20_4,
	input signed [DATA_WIDTH-1:0] in_data_20_5,
	input signed [DATA_WIDTH-1:0] in_data_20_6,
	input signed [DATA_WIDTH-1:0] in_data_20_7,
	input signed [DATA_WIDTH-1:0] in_data_20_8,
	input signed [DATA_WIDTH-1:0] in_data_20_9,
	input signed [DATA_WIDTH-1:0] in_data_20_10,
	input signed [DATA_WIDTH-1:0] in_data_20_11,
	input signed [DATA_WIDTH-1:0] in_data_20_12,
	input signed [DATA_WIDTH-1:0] in_data_20_13,
	input signed [DATA_WIDTH-1:0] in_data_20_14,
	input signed [DATA_WIDTH-1:0] in_data_20_15,
	input signed [DATA_WIDTH-1:0] in_data_20_16,
	input signed [DATA_WIDTH-1:0] in_data_20_17,
	input signed [DATA_WIDTH-1:0] in_data_20_18,
	input signed [DATA_WIDTH-1:0] in_data_20_19,
	input signed [DATA_WIDTH-1:0] in_data_20_20,
	input signed [DATA_WIDTH-1:0] in_data_20_21,
	input signed [DATA_WIDTH-1:0] in_data_20_22,
	input signed [DATA_WIDTH-1:0] in_data_20_23,
	input signed [DATA_WIDTH-1:0] in_data_20_24,
	input signed [DATA_WIDTH-1:0] in_data_20_25,
	input signed [DATA_WIDTH-1:0] in_data_20_26,
	input signed [DATA_WIDTH-1:0] in_data_20_27,
	input signed [DATA_WIDTH-1:0] in_data_20_28,
	input signed [DATA_WIDTH-1:0] in_data_20_29,
	input signed [DATA_WIDTH-1:0] in_data_20_30,
	input signed [DATA_WIDTH-1:0] in_data_20_31,
	input signed [DATA_WIDTH-1:0] in_data_21_0,
	input signed [DATA_WIDTH-1:0] in_data_21_1,
	input signed [DATA_WIDTH-1:0] in_data_21_2,
	input signed [DATA_WIDTH-1:0] in_data_21_3,
	input signed [DATA_WIDTH-1:0] in_data_21_4,
	input signed [DATA_WIDTH-1:0] in_data_21_5,
	input signed [DATA_WIDTH-1:0] in_data_21_6,
	input signed [DATA_WIDTH-1:0] in_data_21_7,
	input signed [DATA_WIDTH-1:0] in_data_21_8,
	input signed [DATA_WIDTH-1:0] in_data_21_9,
	input signed [DATA_WIDTH-1:0] in_data_21_10,
	input signed [DATA_WIDTH-1:0] in_data_21_11,
	input signed [DATA_WIDTH-1:0] in_data_21_12,
	input signed [DATA_WIDTH-1:0] in_data_21_13,
	input signed [DATA_WIDTH-1:0] in_data_21_14,
	input signed [DATA_WIDTH-1:0] in_data_21_15,
	input signed [DATA_WIDTH-1:0] in_data_21_16,
	input signed [DATA_WIDTH-1:0] in_data_21_17,
	input signed [DATA_WIDTH-1:0] in_data_21_18,
	input signed [DATA_WIDTH-1:0] in_data_21_19,
	input signed [DATA_WIDTH-1:0] in_data_21_20,
	input signed [DATA_WIDTH-1:0] in_data_21_21,
	input signed [DATA_WIDTH-1:0] in_data_21_22,
	input signed [DATA_WIDTH-1:0] in_data_21_23,
	input signed [DATA_WIDTH-1:0] in_data_21_24,
	input signed [DATA_WIDTH-1:0] in_data_21_25,
	input signed [DATA_WIDTH-1:0] in_data_21_26,
	input signed [DATA_WIDTH-1:0] in_data_21_27,
	input signed [DATA_WIDTH-1:0] in_data_21_28,
	input signed [DATA_WIDTH-1:0] in_data_21_29,
	input signed [DATA_WIDTH-1:0] in_data_21_30,
	input signed [DATA_WIDTH-1:0] in_data_21_31,
	input signed [DATA_WIDTH-1:0] in_data_22_0,
	input signed [DATA_WIDTH-1:0] in_data_22_1,
	input signed [DATA_WIDTH-1:0] in_data_22_2,
	input signed [DATA_WIDTH-1:0] in_data_22_3,
	input signed [DATA_WIDTH-1:0] in_data_22_4,
	input signed [DATA_WIDTH-1:0] in_data_22_5,
	input signed [DATA_WIDTH-1:0] in_data_22_6,
	input signed [DATA_WIDTH-1:0] in_data_22_7,
	input signed [DATA_WIDTH-1:0] in_data_22_8,
	input signed [DATA_WIDTH-1:0] in_data_22_9,
	input signed [DATA_WIDTH-1:0] in_data_22_10,
	input signed [DATA_WIDTH-1:0] in_data_22_11,
	input signed [DATA_WIDTH-1:0] in_data_22_12,
	input signed [DATA_WIDTH-1:0] in_data_22_13,
	input signed [DATA_WIDTH-1:0] in_data_22_14,
	input signed [DATA_WIDTH-1:0] in_data_22_15,
	input signed [DATA_WIDTH-1:0] in_data_22_16,
	input signed [DATA_WIDTH-1:0] in_data_22_17,
	input signed [DATA_WIDTH-1:0] in_data_22_18,
	input signed [DATA_WIDTH-1:0] in_data_22_19,
	input signed [DATA_WIDTH-1:0] in_data_22_20,
	input signed [DATA_WIDTH-1:0] in_data_22_21,
	input signed [DATA_WIDTH-1:0] in_data_22_22,
	input signed [DATA_WIDTH-1:0] in_data_22_23,
	input signed [DATA_WIDTH-1:0] in_data_22_24,
	input signed [DATA_WIDTH-1:0] in_data_22_25,
	input signed [DATA_WIDTH-1:0] in_data_22_26,
	input signed [DATA_WIDTH-1:0] in_data_22_27,
	input signed [DATA_WIDTH-1:0] in_data_22_28,
	input signed [DATA_WIDTH-1:0] in_data_22_29,
	input signed [DATA_WIDTH-1:0] in_data_22_30,
	input signed [DATA_WIDTH-1:0] in_data_22_31,
	input signed [DATA_WIDTH-1:0] in_data_23_0,
	input signed [DATA_WIDTH-1:0] in_data_23_1,
	input signed [DATA_WIDTH-1:0] in_data_23_2,
	input signed [DATA_WIDTH-1:0] in_data_23_3,
	input signed [DATA_WIDTH-1:0] in_data_23_4,
	input signed [DATA_WIDTH-1:0] in_data_23_5,
	input signed [DATA_WIDTH-1:0] in_data_23_6,
	input signed [DATA_WIDTH-1:0] in_data_23_7,
	input signed [DATA_WIDTH-1:0] in_data_23_8,
	input signed [DATA_WIDTH-1:0] in_data_23_9,
	input signed [DATA_WIDTH-1:0] in_data_23_10,
	input signed [DATA_WIDTH-1:0] in_data_23_11,
	input signed [DATA_WIDTH-1:0] in_data_23_12,
	input signed [DATA_WIDTH-1:0] in_data_23_13,
	input signed [DATA_WIDTH-1:0] in_data_23_14,
	input signed [DATA_WIDTH-1:0] in_data_23_15,
	input signed [DATA_WIDTH-1:0] in_data_23_16,
	input signed [DATA_WIDTH-1:0] in_data_23_17,
	input signed [DATA_WIDTH-1:0] in_data_23_18,
	input signed [DATA_WIDTH-1:0] in_data_23_19,
	input signed [DATA_WIDTH-1:0] in_data_23_20,
	input signed [DATA_WIDTH-1:0] in_data_23_21,
	input signed [DATA_WIDTH-1:0] in_data_23_22,
	input signed [DATA_WIDTH-1:0] in_data_23_23,
	input signed [DATA_WIDTH-1:0] in_data_23_24,
	input signed [DATA_WIDTH-1:0] in_data_23_25,
	input signed [DATA_WIDTH-1:0] in_data_23_26,
	input signed [DATA_WIDTH-1:0] in_data_23_27,
	input signed [DATA_WIDTH-1:0] in_data_23_28,
	input signed [DATA_WIDTH-1:0] in_data_23_29,
	input signed [DATA_WIDTH-1:0] in_data_23_30,
	input signed [DATA_WIDTH-1:0] in_data_23_31,
	input signed [DATA_WIDTH-1:0] in_data_24_0,
	input signed [DATA_WIDTH-1:0] in_data_24_1,
	input signed [DATA_WIDTH-1:0] in_data_24_2,
	input signed [DATA_WIDTH-1:0] in_data_24_3,
	input signed [DATA_WIDTH-1:0] in_data_24_4,
	input signed [DATA_WIDTH-1:0] in_data_24_5,
	input signed [DATA_WIDTH-1:0] in_data_24_6,
	input signed [DATA_WIDTH-1:0] in_data_24_7,
	input signed [DATA_WIDTH-1:0] in_data_24_8,
	input signed [DATA_WIDTH-1:0] in_data_24_9,
	input signed [DATA_WIDTH-1:0] in_data_24_10,
	input signed [DATA_WIDTH-1:0] in_data_24_11,
	input signed [DATA_WIDTH-1:0] in_data_24_12,
	input signed [DATA_WIDTH-1:0] in_data_24_13,
	input signed [DATA_WIDTH-1:0] in_data_24_14,
	input signed [DATA_WIDTH-1:0] in_data_24_15,
	input signed [DATA_WIDTH-1:0] in_data_24_16,
	input signed [DATA_WIDTH-1:0] in_data_24_17,
	input signed [DATA_WIDTH-1:0] in_data_24_18,
	input signed [DATA_WIDTH-1:0] in_data_24_19,
	input signed [DATA_WIDTH-1:0] in_data_24_20,
	input signed [DATA_WIDTH-1:0] in_data_24_21,
	input signed [DATA_WIDTH-1:0] in_data_24_22,
	input signed [DATA_WIDTH-1:0] in_data_24_23,
	input signed [DATA_WIDTH-1:0] in_data_24_24,
	input signed [DATA_WIDTH-1:0] in_data_24_25,
	input signed [DATA_WIDTH-1:0] in_data_24_26,
	input signed [DATA_WIDTH-1:0] in_data_24_27,
	input signed [DATA_WIDTH-1:0] in_data_24_28,
	input signed [DATA_WIDTH-1:0] in_data_24_29,
	input signed [DATA_WIDTH-1:0] in_data_24_30,
	input signed [DATA_WIDTH-1:0] in_data_24_31,
	input signed [DATA_WIDTH-1:0] in_data_25_0,
	input signed [DATA_WIDTH-1:0] in_data_25_1,
	input signed [DATA_WIDTH-1:0] in_data_25_2,
	input signed [DATA_WIDTH-1:0] in_data_25_3,
	input signed [DATA_WIDTH-1:0] in_data_25_4,
	input signed [DATA_WIDTH-1:0] in_data_25_5,
	input signed [DATA_WIDTH-1:0] in_data_25_6,
	input signed [DATA_WIDTH-1:0] in_data_25_7,
	input signed [DATA_WIDTH-1:0] in_data_25_8,
	input signed [DATA_WIDTH-1:0] in_data_25_9,
	input signed [DATA_WIDTH-1:0] in_data_25_10,
	input signed [DATA_WIDTH-1:0] in_data_25_11,
	input signed [DATA_WIDTH-1:0] in_data_25_12,
	input signed [DATA_WIDTH-1:0] in_data_25_13,
	input signed [DATA_WIDTH-1:0] in_data_25_14,
	input signed [DATA_WIDTH-1:0] in_data_25_15,
	input signed [DATA_WIDTH-1:0] in_data_25_16,
	input signed [DATA_WIDTH-1:0] in_data_25_17,
	input signed [DATA_WIDTH-1:0] in_data_25_18,
	input signed [DATA_WIDTH-1:0] in_data_25_19,
	input signed [DATA_WIDTH-1:0] in_data_25_20,
	input signed [DATA_WIDTH-1:0] in_data_25_21,
	input signed [DATA_WIDTH-1:0] in_data_25_22,
	input signed [DATA_WIDTH-1:0] in_data_25_23,
	input signed [DATA_WIDTH-1:0] in_data_25_24,
	input signed [DATA_WIDTH-1:0] in_data_25_25,
	input signed [DATA_WIDTH-1:0] in_data_25_26,
	input signed [DATA_WIDTH-1:0] in_data_25_27,
	input signed [DATA_WIDTH-1:0] in_data_25_28,
	input signed [DATA_WIDTH-1:0] in_data_25_29,
	input signed [DATA_WIDTH-1:0] in_data_25_30,
	input signed [DATA_WIDTH-1:0] in_data_25_31,
	input signed [DATA_WIDTH-1:0] in_data_26_0,
	input signed [DATA_WIDTH-1:0] in_data_26_1,
	input signed [DATA_WIDTH-1:0] in_data_26_2,
	input signed [DATA_WIDTH-1:0] in_data_26_3,
	input signed [DATA_WIDTH-1:0] in_data_26_4,
	input signed [DATA_WIDTH-1:0] in_data_26_5,
	input signed [DATA_WIDTH-1:0] in_data_26_6,
	input signed [DATA_WIDTH-1:0] in_data_26_7,
	input signed [DATA_WIDTH-1:0] in_data_26_8,
	input signed [DATA_WIDTH-1:0] in_data_26_9,
	input signed [DATA_WIDTH-1:0] in_data_26_10,
	input signed [DATA_WIDTH-1:0] in_data_26_11,
	input signed [DATA_WIDTH-1:0] in_data_26_12,
	input signed [DATA_WIDTH-1:0] in_data_26_13,
	input signed [DATA_WIDTH-1:0] in_data_26_14,
	input signed [DATA_WIDTH-1:0] in_data_26_15,
	input signed [DATA_WIDTH-1:0] in_data_26_16,
	input signed [DATA_WIDTH-1:0] in_data_26_17,
	input signed [DATA_WIDTH-1:0] in_data_26_18,
	input signed [DATA_WIDTH-1:0] in_data_26_19,
	input signed [DATA_WIDTH-1:0] in_data_26_20,
	input signed [DATA_WIDTH-1:0] in_data_26_21,
	input signed [DATA_WIDTH-1:0] in_data_26_22,
	input signed [DATA_WIDTH-1:0] in_data_26_23,
	input signed [DATA_WIDTH-1:0] in_data_26_24,
	input signed [DATA_WIDTH-1:0] in_data_26_25,
	input signed [DATA_WIDTH-1:0] in_data_26_26,
	input signed [DATA_WIDTH-1:0] in_data_26_27,
	input signed [DATA_WIDTH-1:0] in_data_26_28,
	input signed [DATA_WIDTH-1:0] in_data_26_29,
	input signed [DATA_WIDTH-1:0] in_data_26_30,
	input signed [DATA_WIDTH-1:0] in_data_26_31,
	input signed [DATA_WIDTH-1:0] in_data_27_0,
	input signed [DATA_WIDTH-1:0] in_data_27_1,
	input signed [DATA_WIDTH-1:0] in_data_27_2,
	input signed [DATA_WIDTH-1:0] in_data_27_3,
	input signed [DATA_WIDTH-1:0] in_data_27_4,
	input signed [DATA_WIDTH-1:0] in_data_27_5,
	input signed [DATA_WIDTH-1:0] in_data_27_6,
	input signed [DATA_WIDTH-1:0] in_data_27_7,
	input signed [DATA_WIDTH-1:0] in_data_27_8,
	input signed [DATA_WIDTH-1:0] in_data_27_9,
	input signed [DATA_WIDTH-1:0] in_data_27_10,
	input signed [DATA_WIDTH-1:0] in_data_27_11,
	input signed [DATA_WIDTH-1:0] in_data_27_12,
	input signed [DATA_WIDTH-1:0] in_data_27_13,
	input signed [DATA_WIDTH-1:0] in_data_27_14,
	input signed [DATA_WIDTH-1:0] in_data_27_15,
	input signed [DATA_WIDTH-1:0] in_data_27_16,
	input signed [DATA_WIDTH-1:0] in_data_27_17,
	input signed [DATA_WIDTH-1:0] in_data_27_18,
	input signed [DATA_WIDTH-1:0] in_data_27_19,
	input signed [DATA_WIDTH-1:0] in_data_27_20,
	input signed [DATA_WIDTH-1:0] in_data_27_21,
	input signed [DATA_WIDTH-1:0] in_data_27_22,
	input signed [DATA_WIDTH-1:0] in_data_27_23,
	input signed [DATA_WIDTH-1:0] in_data_27_24,
	input signed [DATA_WIDTH-1:0] in_data_27_25,
	input signed [DATA_WIDTH-1:0] in_data_27_26,
	input signed [DATA_WIDTH-1:0] in_data_27_27,
	input signed [DATA_WIDTH-1:0] in_data_27_28,
	input signed [DATA_WIDTH-1:0] in_data_27_29,
	input signed [DATA_WIDTH-1:0] in_data_27_30,
	input signed [DATA_WIDTH-1:0] in_data_27_31,
	input signed [DATA_WIDTH-1:0] in_data_28_0,
	input signed [DATA_WIDTH-1:0] in_data_28_1,
	input signed [DATA_WIDTH-1:0] in_data_28_2,
	input signed [DATA_WIDTH-1:0] in_data_28_3,
	input signed [DATA_WIDTH-1:0] in_data_28_4,
	input signed [DATA_WIDTH-1:0] in_data_28_5,
	input signed [DATA_WIDTH-1:0] in_data_28_6,
	input signed [DATA_WIDTH-1:0] in_data_28_7,
	input signed [DATA_WIDTH-1:0] in_data_28_8,
	input signed [DATA_WIDTH-1:0] in_data_28_9,
	input signed [DATA_WIDTH-1:0] in_data_28_10,
	input signed [DATA_WIDTH-1:0] in_data_28_11,
	input signed [DATA_WIDTH-1:0] in_data_28_12,
	input signed [DATA_WIDTH-1:0] in_data_28_13,
	input signed [DATA_WIDTH-1:0] in_data_28_14,
	input signed [DATA_WIDTH-1:0] in_data_28_15,
	input signed [DATA_WIDTH-1:0] in_data_28_16,
	input signed [DATA_WIDTH-1:0] in_data_28_17,
	input signed [DATA_WIDTH-1:0] in_data_28_18,
	input signed [DATA_WIDTH-1:0] in_data_28_19,
	input signed [DATA_WIDTH-1:0] in_data_28_20,
	input signed [DATA_WIDTH-1:0] in_data_28_21,
	input signed [DATA_WIDTH-1:0] in_data_28_22,
	input signed [DATA_WIDTH-1:0] in_data_28_23,
	input signed [DATA_WIDTH-1:0] in_data_28_24,
	input signed [DATA_WIDTH-1:0] in_data_28_25,
	input signed [DATA_WIDTH-1:0] in_data_28_26,
	input signed [DATA_WIDTH-1:0] in_data_28_27,
	input signed [DATA_WIDTH-1:0] in_data_28_28,
	input signed [DATA_WIDTH-1:0] in_data_28_29,
	input signed [DATA_WIDTH-1:0] in_data_28_30,
	input signed [DATA_WIDTH-1:0] in_data_28_31,
	input signed [DATA_WIDTH-1:0] in_data_29_0,
	input signed [DATA_WIDTH-1:0] in_data_29_1,
	input signed [DATA_WIDTH-1:0] in_data_29_2,
	input signed [DATA_WIDTH-1:0] in_data_29_3,
	input signed [DATA_WIDTH-1:0] in_data_29_4,
	input signed [DATA_WIDTH-1:0] in_data_29_5,
	input signed [DATA_WIDTH-1:0] in_data_29_6,
	input signed [DATA_WIDTH-1:0] in_data_29_7,
	input signed [DATA_WIDTH-1:0] in_data_29_8,
	input signed [DATA_WIDTH-1:0] in_data_29_9,
	input signed [DATA_WIDTH-1:0] in_data_29_10,
	input signed [DATA_WIDTH-1:0] in_data_29_11,
	input signed [DATA_WIDTH-1:0] in_data_29_12,
	input signed [DATA_WIDTH-1:0] in_data_29_13,
	input signed [DATA_WIDTH-1:0] in_data_29_14,
	input signed [DATA_WIDTH-1:0] in_data_29_15,
	input signed [DATA_WIDTH-1:0] in_data_29_16,
	input signed [DATA_WIDTH-1:0] in_data_29_17,
	input signed [DATA_WIDTH-1:0] in_data_29_18,
	input signed [DATA_WIDTH-1:0] in_data_29_19,
	input signed [DATA_WIDTH-1:0] in_data_29_20,
	input signed [DATA_WIDTH-1:0] in_data_29_21,
	input signed [DATA_WIDTH-1:0] in_data_29_22,
	input signed [DATA_WIDTH-1:0] in_data_29_23,
	input signed [DATA_WIDTH-1:0] in_data_29_24,
	input signed [DATA_WIDTH-1:0] in_data_29_25,
	input signed [DATA_WIDTH-1:0] in_data_29_26,
	input signed [DATA_WIDTH-1:0] in_data_29_27,
	input signed [DATA_WIDTH-1:0] in_data_29_28,
	input signed [DATA_WIDTH-1:0] in_data_29_29,
	input signed [DATA_WIDTH-1:0] in_data_29_30,
	input signed [DATA_WIDTH-1:0] in_data_29_31,
	input signed [DATA_WIDTH-1:0] in_data_30_0,
	input signed [DATA_WIDTH-1:0] in_data_30_1,
	input signed [DATA_WIDTH-1:0] in_data_30_2,
	input signed [DATA_WIDTH-1:0] in_data_30_3,
	input signed [DATA_WIDTH-1:0] in_data_30_4,
	input signed [DATA_WIDTH-1:0] in_data_30_5,
	input signed [DATA_WIDTH-1:0] in_data_30_6,
	input signed [DATA_WIDTH-1:0] in_data_30_7,
	input signed [DATA_WIDTH-1:0] in_data_30_8,
	input signed [DATA_WIDTH-1:0] in_data_30_9,
	input signed [DATA_WIDTH-1:0] in_data_30_10,
	input signed [DATA_WIDTH-1:0] in_data_30_11,
	input signed [DATA_WIDTH-1:0] in_data_30_12,
	input signed [DATA_WIDTH-1:0] in_data_30_13,
	input signed [DATA_WIDTH-1:0] in_data_30_14,
	input signed [DATA_WIDTH-1:0] in_data_30_15,
	input signed [DATA_WIDTH-1:0] in_data_30_16,
	input signed [DATA_WIDTH-1:0] in_data_30_17,
	input signed [DATA_WIDTH-1:0] in_data_30_18,
	input signed [DATA_WIDTH-1:0] in_data_30_19,
	input signed [DATA_WIDTH-1:0] in_data_30_20,
	input signed [DATA_WIDTH-1:0] in_data_30_21,
	input signed [DATA_WIDTH-1:0] in_data_30_22,
	input signed [DATA_WIDTH-1:0] in_data_30_23,
	input signed [DATA_WIDTH-1:0] in_data_30_24,
	input signed [DATA_WIDTH-1:0] in_data_30_25,
	input signed [DATA_WIDTH-1:0] in_data_30_26,
	input signed [DATA_WIDTH-1:0] in_data_30_27,
	input signed [DATA_WIDTH-1:0] in_data_30_28,
	input signed [DATA_WIDTH-1:0] in_data_30_29,
	input signed [DATA_WIDTH-1:0] in_data_30_30,
	input signed [DATA_WIDTH-1:0] in_data_30_31,
	input signed [DATA_WIDTH-1:0] in_data_31_0,
	input signed [DATA_WIDTH-1:0] in_data_31_1,
	input signed [DATA_WIDTH-1:0] in_data_31_2,
	input signed [DATA_WIDTH-1:0] in_data_31_3,
	input signed [DATA_WIDTH-1:0] in_data_31_4,
	input signed [DATA_WIDTH-1:0] in_data_31_5,
	input signed [DATA_WIDTH-1:0] in_data_31_6,
	input signed [DATA_WIDTH-1:0] in_data_31_7,
	input signed [DATA_WIDTH-1:0] in_data_31_8,
	input signed [DATA_WIDTH-1:0] in_data_31_9,
	input signed [DATA_WIDTH-1:0] in_data_31_10,
	input signed [DATA_WIDTH-1:0] in_data_31_11,
	input signed [DATA_WIDTH-1:0] in_data_31_12,
	input signed [DATA_WIDTH-1:0] in_data_31_13,
	input signed [DATA_WIDTH-1:0] in_data_31_14,
	input signed [DATA_WIDTH-1:0] in_data_31_15,
	input signed [DATA_WIDTH-1:0] in_data_31_16,
	input signed [DATA_WIDTH-1:0] in_data_31_17,
	input signed [DATA_WIDTH-1:0] in_data_31_18,
	input signed [DATA_WIDTH-1:0] in_data_31_19,
	input signed [DATA_WIDTH-1:0] in_data_31_20,
	input signed [DATA_WIDTH-1:0] in_data_31_21,
	input signed [DATA_WIDTH-1:0] in_data_31_22,
	input signed [DATA_WIDTH-1:0] in_data_31_23,
	input signed [DATA_WIDTH-1:0] in_data_31_24,
	input signed [DATA_WIDTH-1:0] in_data_31_25,
	input signed [DATA_WIDTH-1:0] in_data_31_26,
	input signed [DATA_WIDTH-1:0] in_data_31_27,
	input signed [DATA_WIDTH-1:0] in_data_31_28,
	input signed [DATA_WIDTH-1:0] in_data_31_29,
	input signed [DATA_WIDTH-1:0] in_data_31_30,
	input signed [DATA_WIDTH-1:0] in_data_31_31,
	output reg signed [DATA_WIDTH-1:0] out_data
);

  // Perform mux operation
  always @ (select) begin
    case (select)
			10'b0000000000 : out_data <= in_data_0_0;
			10'b0000000001 : out_data <= in_data_0_1;
			10'b0000000010 : out_data <= in_data_0_2;
			10'b0000000011 : out_data <= in_data_0_3;
			10'b0000000100 : out_data <= in_data_0_4;
			10'b0000000101 : out_data <= in_data_0_5;
			10'b0000000110 : out_data <= in_data_0_6;
			10'b0000000111 : out_data <= in_data_0_7;
			10'b0000001000 : out_data <= in_data_0_8;
			10'b0000001001 : out_data <= in_data_0_9;
			10'b0000001010 : out_data <= in_data_0_10;
			10'b0000001011 : out_data <= in_data_0_11;
			10'b0000001100 : out_data <= in_data_0_12;
			10'b0000001101 : out_data <= in_data_0_13;
			10'b0000001110 : out_data <= in_data_0_14;
			10'b0000001111 : out_data <= in_data_0_15;
			10'b0000010000 : out_data <= in_data_0_16;
			10'b0000010001 : out_data <= in_data_0_17;
			10'b0000010010 : out_data <= in_data_0_18;
			10'b0000010011 : out_data <= in_data_0_19;
			10'b0000010100 : out_data <= in_data_0_20;
			10'b0000010101 : out_data <= in_data_0_21;
			10'b0000010110 : out_data <= in_data_0_22;
			10'b0000010111 : out_data <= in_data_0_23;
			10'b0000011000 : out_data <= in_data_0_24;
			10'b0000011001 : out_data <= in_data_0_25;
			10'b0000011010 : out_data <= in_data_0_26;
			10'b0000011011 : out_data <= in_data_0_27;
			10'b0000011100 : out_data <= in_data_0_28;
			10'b0000011101 : out_data <= in_data_0_29;
			10'b0000011110 : out_data <= in_data_0_30;
			10'b0000011111 : out_data <= in_data_0_31;
			10'b0000100000 : out_data <= in_data_1_0;
			10'b0000100001 : out_data <= in_data_1_1;
			10'b0000100010 : out_data <= in_data_1_2;
			10'b0000100011 : out_data <= in_data_1_3;
			10'b0000100100 : out_data <= in_data_1_4;
			10'b0000100101 : out_data <= in_data_1_5;
			10'b0000100110 : out_data <= in_data_1_6;
			10'b0000100111 : out_data <= in_data_1_7;
			10'b0000101000 : out_data <= in_data_1_8;
			10'b0000101001 : out_data <= in_data_1_9;
			10'b0000101010 : out_data <= in_data_1_10;
			10'b0000101011 : out_data <= in_data_1_11;
			10'b0000101100 : out_data <= in_data_1_12;
			10'b0000101101 : out_data <= in_data_1_13;
			10'b0000101110 : out_data <= in_data_1_14;
			10'b0000101111 : out_data <= in_data_1_15;
			10'b0000110000 : out_data <= in_data_1_16;
			10'b0000110001 : out_data <= in_data_1_17;
			10'b0000110010 : out_data <= in_data_1_18;
			10'b0000110011 : out_data <= in_data_1_19;
			10'b0000110100 : out_data <= in_data_1_20;
			10'b0000110101 : out_data <= in_data_1_21;
			10'b0000110110 : out_data <= in_data_1_22;
			10'b0000110111 : out_data <= in_data_1_23;
			10'b0000111000 : out_data <= in_data_1_24;
			10'b0000111001 : out_data <= in_data_1_25;
			10'b0000111010 : out_data <= in_data_1_26;
			10'b0000111011 : out_data <= in_data_1_27;
			10'b0000111100 : out_data <= in_data_1_28;
			10'b0000111101 : out_data <= in_data_1_29;
			10'b0000111110 : out_data <= in_data_1_30;
			10'b0000111111 : out_data <= in_data_1_31;
			10'b0001000000 : out_data <= in_data_2_0;
			10'b0001000001 : out_data <= in_data_2_1;
			10'b0001000010 : out_data <= in_data_2_2;
			10'b0001000011 : out_data <= in_data_2_3;
			10'b0001000100 : out_data <= in_data_2_4;
			10'b0001000101 : out_data <= in_data_2_5;
			10'b0001000110 : out_data <= in_data_2_6;
			10'b0001000111 : out_data <= in_data_2_7;
			10'b0001001000 : out_data <= in_data_2_8;
			10'b0001001001 : out_data <= in_data_2_9;
			10'b0001001010 : out_data <= in_data_2_10;
			10'b0001001011 : out_data <= in_data_2_11;
			10'b0001001100 : out_data <= in_data_2_12;
			10'b0001001101 : out_data <= in_data_2_13;
			10'b0001001110 : out_data <= in_data_2_14;
			10'b0001001111 : out_data <= in_data_2_15;
			10'b0001010000 : out_data <= in_data_2_16;
			10'b0001010001 : out_data <= in_data_2_17;
			10'b0001010010 : out_data <= in_data_2_18;
			10'b0001010011 : out_data <= in_data_2_19;
			10'b0001010100 : out_data <= in_data_2_20;
			10'b0001010101 : out_data <= in_data_2_21;
			10'b0001010110 : out_data <= in_data_2_22;
			10'b0001010111 : out_data <= in_data_2_23;
			10'b0001011000 : out_data <= in_data_2_24;
			10'b0001011001 : out_data <= in_data_2_25;
			10'b0001011010 : out_data <= in_data_2_26;
			10'b0001011011 : out_data <= in_data_2_27;
			10'b0001011100 : out_data <= in_data_2_28;
			10'b0001011101 : out_data <= in_data_2_29;
			10'b0001011110 : out_data <= in_data_2_30;
			10'b0001011111 : out_data <= in_data_2_31;
			10'b0001100000 : out_data <= in_data_3_0;
			10'b0001100001 : out_data <= in_data_3_1;
			10'b0001100010 : out_data <= in_data_3_2;
			10'b0001100011 : out_data <= in_data_3_3;
			10'b0001100100 : out_data <= in_data_3_4;
			10'b0001100101 : out_data <= in_data_3_5;
			10'b0001100110 : out_data <= in_data_3_6;
			10'b0001100111 : out_data <= in_data_3_7;
			10'b0001101000 : out_data <= in_data_3_8;
			10'b0001101001 : out_data <= in_data_3_9;
			10'b0001101010 : out_data <= in_data_3_10;
			10'b0001101011 : out_data <= in_data_3_11;
			10'b0001101100 : out_data <= in_data_3_12;
			10'b0001101101 : out_data <= in_data_3_13;
			10'b0001101110 : out_data <= in_data_3_14;
			10'b0001101111 : out_data <= in_data_3_15;
			10'b0001110000 : out_data <= in_data_3_16;
			10'b0001110001 : out_data <= in_data_3_17;
			10'b0001110010 : out_data <= in_data_3_18;
			10'b0001110011 : out_data <= in_data_3_19;
			10'b0001110100 : out_data <= in_data_3_20;
			10'b0001110101 : out_data <= in_data_3_21;
			10'b0001110110 : out_data <= in_data_3_22;
			10'b0001110111 : out_data <= in_data_3_23;
			10'b0001111000 : out_data <= in_data_3_24;
			10'b0001111001 : out_data <= in_data_3_25;
			10'b0001111010 : out_data <= in_data_3_26;
			10'b0001111011 : out_data <= in_data_3_27;
			10'b0001111100 : out_data <= in_data_3_28;
			10'b0001111101 : out_data <= in_data_3_29;
			10'b0001111110 : out_data <= in_data_3_30;
			10'b0001111111 : out_data <= in_data_3_31;
			10'b0010000000 : out_data <= in_data_4_0;
			10'b0010000001 : out_data <= in_data_4_1;
			10'b0010000010 : out_data <= in_data_4_2;
			10'b0010000011 : out_data <= in_data_4_3;
			10'b0010000100 : out_data <= in_data_4_4;
			10'b0010000101 : out_data <= in_data_4_5;
			10'b0010000110 : out_data <= in_data_4_6;
			10'b0010000111 : out_data <= in_data_4_7;
			10'b0010001000 : out_data <= in_data_4_8;
			10'b0010001001 : out_data <= in_data_4_9;
			10'b0010001010 : out_data <= in_data_4_10;
			10'b0010001011 : out_data <= in_data_4_11;
			10'b0010001100 : out_data <= in_data_4_12;
			10'b0010001101 : out_data <= in_data_4_13;
			10'b0010001110 : out_data <= in_data_4_14;
			10'b0010001111 : out_data <= in_data_4_15;
			10'b0010010000 : out_data <= in_data_4_16;
			10'b0010010001 : out_data <= in_data_4_17;
			10'b0010010010 : out_data <= in_data_4_18;
			10'b0010010011 : out_data <= in_data_4_19;
			10'b0010010100 : out_data <= in_data_4_20;
			10'b0010010101 : out_data <= in_data_4_21;
			10'b0010010110 : out_data <= in_data_4_22;
			10'b0010010111 : out_data <= in_data_4_23;
			10'b0010011000 : out_data <= in_data_4_24;
			10'b0010011001 : out_data <= in_data_4_25;
			10'b0010011010 : out_data <= in_data_4_26;
			10'b0010011011 : out_data <= in_data_4_27;
			10'b0010011100 : out_data <= in_data_4_28;
			10'b0010011101 : out_data <= in_data_4_29;
			10'b0010011110 : out_data <= in_data_4_30;
			10'b0010011111 : out_data <= in_data_4_31;
			10'b0010100000 : out_data <= in_data_5_0;
			10'b0010100001 : out_data <= in_data_5_1;
			10'b0010100010 : out_data <= in_data_5_2;
			10'b0010100011 : out_data <= in_data_5_3;
			10'b0010100100 : out_data <= in_data_5_4;
			10'b0010100101 : out_data <= in_data_5_5;
			10'b0010100110 : out_data <= in_data_5_6;
			10'b0010100111 : out_data <= in_data_5_7;
			10'b0010101000 : out_data <= in_data_5_8;
			10'b0010101001 : out_data <= in_data_5_9;
			10'b0010101010 : out_data <= in_data_5_10;
			10'b0010101011 : out_data <= in_data_5_11;
			10'b0010101100 : out_data <= in_data_5_12;
			10'b0010101101 : out_data <= in_data_5_13;
			10'b0010101110 : out_data <= in_data_5_14;
			10'b0010101111 : out_data <= in_data_5_15;
			10'b0010110000 : out_data <= in_data_5_16;
			10'b0010110001 : out_data <= in_data_5_17;
			10'b0010110010 : out_data <= in_data_5_18;
			10'b0010110011 : out_data <= in_data_5_19;
			10'b0010110100 : out_data <= in_data_5_20;
			10'b0010110101 : out_data <= in_data_5_21;
			10'b0010110110 : out_data <= in_data_5_22;
			10'b0010110111 : out_data <= in_data_5_23;
			10'b0010111000 : out_data <= in_data_5_24;
			10'b0010111001 : out_data <= in_data_5_25;
			10'b0010111010 : out_data <= in_data_5_26;
			10'b0010111011 : out_data <= in_data_5_27;
			10'b0010111100 : out_data <= in_data_5_28;
			10'b0010111101 : out_data <= in_data_5_29;
			10'b0010111110 : out_data <= in_data_5_30;
			10'b0010111111 : out_data <= in_data_5_31;
			10'b0011000000 : out_data <= in_data_6_0;
			10'b0011000001 : out_data <= in_data_6_1;
			10'b0011000010 : out_data <= in_data_6_2;
			10'b0011000011 : out_data <= in_data_6_3;
			10'b0011000100 : out_data <= in_data_6_4;
			10'b0011000101 : out_data <= in_data_6_5;
			10'b0011000110 : out_data <= in_data_6_6;
			10'b0011000111 : out_data <= in_data_6_7;
			10'b0011001000 : out_data <= in_data_6_8;
			10'b0011001001 : out_data <= in_data_6_9;
			10'b0011001010 : out_data <= in_data_6_10;
			10'b0011001011 : out_data <= in_data_6_11;
			10'b0011001100 : out_data <= in_data_6_12;
			10'b0011001101 : out_data <= in_data_6_13;
			10'b0011001110 : out_data <= in_data_6_14;
			10'b0011001111 : out_data <= in_data_6_15;
			10'b0011010000 : out_data <= in_data_6_16;
			10'b0011010001 : out_data <= in_data_6_17;
			10'b0011010010 : out_data <= in_data_6_18;
			10'b0011010011 : out_data <= in_data_6_19;
			10'b0011010100 : out_data <= in_data_6_20;
			10'b0011010101 : out_data <= in_data_6_21;
			10'b0011010110 : out_data <= in_data_6_22;
			10'b0011010111 : out_data <= in_data_6_23;
			10'b0011011000 : out_data <= in_data_6_24;
			10'b0011011001 : out_data <= in_data_6_25;
			10'b0011011010 : out_data <= in_data_6_26;
			10'b0011011011 : out_data <= in_data_6_27;
			10'b0011011100 : out_data <= in_data_6_28;
			10'b0011011101 : out_data <= in_data_6_29;
			10'b0011011110 : out_data <= in_data_6_30;
			10'b0011011111 : out_data <= in_data_6_31;
			10'b0011100000 : out_data <= in_data_7_0;
			10'b0011100001 : out_data <= in_data_7_1;
			10'b0011100010 : out_data <= in_data_7_2;
			10'b0011100011 : out_data <= in_data_7_3;
			10'b0011100100 : out_data <= in_data_7_4;
			10'b0011100101 : out_data <= in_data_7_5;
			10'b0011100110 : out_data <= in_data_7_6;
			10'b0011100111 : out_data <= in_data_7_7;
			10'b0011101000 : out_data <= in_data_7_8;
			10'b0011101001 : out_data <= in_data_7_9;
			10'b0011101010 : out_data <= in_data_7_10;
			10'b0011101011 : out_data <= in_data_7_11;
			10'b0011101100 : out_data <= in_data_7_12;
			10'b0011101101 : out_data <= in_data_7_13;
			10'b0011101110 : out_data <= in_data_7_14;
			10'b0011101111 : out_data <= in_data_7_15;
			10'b0011110000 : out_data <= in_data_7_16;
			10'b0011110001 : out_data <= in_data_7_17;
			10'b0011110010 : out_data <= in_data_7_18;
			10'b0011110011 : out_data <= in_data_7_19;
			10'b0011110100 : out_data <= in_data_7_20;
			10'b0011110101 : out_data <= in_data_7_21;
			10'b0011110110 : out_data <= in_data_7_22;
			10'b0011110111 : out_data <= in_data_7_23;
			10'b0011111000 : out_data <= in_data_7_24;
			10'b0011111001 : out_data <= in_data_7_25;
			10'b0011111010 : out_data <= in_data_7_26;
			10'b0011111011 : out_data <= in_data_7_27;
			10'b0011111100 : out_data <= in_data_7_28;
			10'b0011111101 : out_data <= in_data_7_29;
			10'b0011111110 : out_data <= in_data_7_30;
			10'b0011111111 : out_data <= in_data_7_31;
			10'b0100000000 : out_data <= in_data_8_0;
			10'b0100000001 : out_data <= in_data_8_1;
			10'b0100000010 : out_data <= in_data_8_2;
			10'b0100000011 : out_data <= in_data_8_3;
			10'b0100000100 : out_data <= in_data_8_4;
			10'b0100000101 : out_data <= in_data_8_5;
			10'b0100000110 : out_data <= in_data_8_6;
			10'b0100000111 : out_data <= in_data_8_7;
			10'b0100001000 : out_data <= in_data_8_8;
			10'b0100001001 : out_data <= in_data_8_9;
			10'b0100001010 : out_data <= in_data_8_10;
			10'b0100001011 : out_data <= in_data_8_11;
			10'b0100001100 : out_data <= in_data_8_12;
			10'b0100001101 : out_data <= in_data_8_13;
			10'b0100001110 : out_data <= in_data_8_14;
			10'b0100001111 : out_data <= in_data_8_15;
			10'b0100010000 : out_data <= in_data_8_16;
			10'b0100010001 : out_data <= in_data_8_17;
			10'b0100010010 : out_data <= in_data_8_18;
			10'b0100010011 : out_data <= in_data_8_19;
			10'b0100010100 : out_data <= in_data_8_20;
			10'b0100010101 : out_data <= in_data_8_21;
			10'b0100010110 : out_data <= in_data_8_22;
			10'b0100010111 : out_data <= in_data_8_23;
			10'b0100011000 : out_data <= in_data_8_24;
			10'b0100011001 : out_data <= in_data_8_25;
			10'b0100011010 : out_data <= in_data_8_26;
			10'b0100011011 : out_data <= in_data_8_27;
			10'b0100011100 : out_data <= in_data_8_28;
			10'b0100011101 : out_data <= in_data_8_29;
			10'b0100011110 : out_data <= in_data_8_30;
			10'b0100011111 : out_data <= in_data_8_31;
			10'b0100100000 : out_data <= in_data_9_0;
			10'b0100100001 : out_data <= in_data_9_1;
			10'b0100100010 : out_data <= in_data_9_2;
			10'b0100100011 : out_data <= in_data_9_3;
			10'b0100100100 : out_data <= in_data_9_4;
			10'b0100100101 : out_data <= in_data_9_5;
			10'b0100100110 : out_data <= in_data_9_6;
			10'b0100100111 : out_data <= in_data_9_7;
			10'b0100101000 : out_data <= in_data_9_8;
			10'b0100101001 : out_data <= in_data_9_9;
			10'b0100101010 : out_data <= in_data_9_10;
			10'b0100101011 : out_data <= in_data_9_11;
			10'b0100101100 : out_data <= in_data_9_12;
			10'b0100101101 : out_data <= in_data_9_13;
			10'b0100101110 : out_data <= in_data_9_14;
			10'b0100101111 : out_data <= in_data_9_15;
			10'b0100110000 : out_data <= in_data_9_16;
			10'b0100110001 : out_data <= in_data_9_17;
			10'b0100110010 : out_data <= in_data_9_18;
			10'b0100110011 : out_data <= in_data_9_19;
			10'b0100110100 : out_data <= in_data_9_20;
			10'b0100110101 : out_data <= in_data_9_21;
			10'b0100110110 : out_data <= in_data_9_22;
			10'b0100110111 : out_data <= in_data_9_23;
			10'b0100111000 : out_data <= in_data_9_24;
			10'b0100111001 : out_data <= in_data_9_25;
			10'b0100111010 : out_data <= in_data_9_26;
			10'b0100111011 : out_data <= in_data_9_27;
			10'b0100111100 : out_data <= in_data_9_28;
			10'b0100111101 : out_data <= in_data_9_29;
			10'b0100111110 : out_data <= in_data_9_30;
			10'b0100111111 : out_data <= in_data_9_31;
			10'b0101000000 : out_data <= in_data_10_0;
			10'b0101000001 : out_data <= in_data_10_1;
			10'b0101000010 : out_data <= in_data_10_2;
			10'b0101000011 : out_data <= in_data_10_3;
			10'b0101000100 : out_data <= in_data_10_4;
			10'b0101000101 : out_data <= in_data_10_5;
			10'b0101000110 : out_data <= in_data_10_6;
			10'b0101000111 : out_data <= in_data_10_7;
			10'b0101001000 : out_data <= in_data_10_8;
			10'b0101001001 : out_data <= in_data_10_9;
			10'b0101001010 : out_data <= in_data_10_10;
			10'b0101001011 : out_data <= in_data_10_11;
			10'b0101001100 : out_data <= in_data_10_12;
			10'b0101001101 : out_data <= in_data_10_13;
			10'b0101001110 : out_data <= in_data_10_14;
			10'b0101001111 : out_data <= in_data_10_15;
			10'b0101010000 : out_data <= in_data_10_16;
			10'b0101010001 : out_data <= in_data_10_17;
			10'b0101010010 : out_data <= in_data_10_18;
			10'b0101010011 : out_data <= in_data_10_19;
			10'b0101010100 : out_data <= in_data_10_20;
			10'b0101010101 : out_data <= in_data_10_21;
			10'b0101010110 : out_data <= in_data_10_22;
			10'b0101010111 : out_data <= in_data_10_23;
			10'b0101011000 : out_data <= in_data_10_24;
			10'b0101011001 : out_data <= in_data_10_25;
			10'b0101011010 : out_data <= in_data_10_26;
			10'b0101011011 : out_data <= in_data_10_27;
			10'b0101011100 : out_data <= in_data_10_28;
			10'b0101011101 : out_data <= in_data_10_29;
			10'b0101011110 : out_data <= in_data_10_30;
			10'b0101011111 : out_data <= in_data_10_31;
			10'b0101100000 : out_data <= in_data_11_0;
			10'b0101100001 : out_data <= in_data_11_1;
			10'b0101100010 : out_data <= in_data_11_2;
			10'b0101100011 : out_data <= in_data_11_3;
			10'b0101100100 : out_data <= in_data_11_4;
			10'b0101100101 : out_data <= in_data_11_5;
			10'b0101100110 : out_data <= in_data_11_6;
			10'b0101100111 : out_data <= in_data_11_7;
			10'b0101101000 : out_data <= in_data_11_8;
			10'b0101101001 : out_data <= in_data_11_9;
			10'b0101101010 : out_data <= in_data_11_10;
			10'b0101101011 : out_data <= in_data_11_11;
			10'b0101101100 : out_data <= in_data_11_12;
			10'b0101101101 : out_data <= in_data_11_13;
			10'b0101101110 : out_data <= in_data_11_14;
			10'b0101101111 : out_data <= in_data_11_15;
			10'b0101110000 : out_data <= in_data_11_16;
			10'b0101110001 : out_data <= in_data_11_17;
			10'b0101110010 : out_data <= in_data_11_18;
			10'b0101110011 : out_data <= in_data_11_19;
			10'b0101110100 : out_data <= in_data_11_20;
			10'b0101110101 : out_data <= in_data_11_21;
			10'b0101110110 : out_data <= in_data_11_22;
			10'b0101110111 : out_data <= in_data_11_23;
			10'b0101111000 : out_data <= in_data_11_24;
			10'b0101111001 : out_data <= in_data_11_25;
			10'b0101111010 : out_data <= in_data_11_26;
			10'b0101111011 : out_data <= in_data_11_27;
			10'b0101111100 : out_data <= in_data_11_28;
			10'b0101111101 : out_data <= in_data_11_29;
			10'b0101111110 : out_data <= in_data_11_30;
			10'b0101111111 : out_data <= in_data_11_31;
			10'b0110000000 : out_data <= in_data_12_0;
			10'b0110000001 : out_data <= in_data_12_1;
			10'b0110000010 : out_data <= in_data_12_2;
			10'b0110000011 : out_data <= in_data_12_3;
			10'b0110000100 : out_data <= in_data_12_4;
			10'b0110000101 : out_data <= in_data_12_5;
			10'b0110000110 : out_data <= in_data_12_6;
			10'b0110000111 : out_data <= in_data_12_7;
			10'b0110001000 : out_data <= in_data_12_8;
			10'b0110001001 : out_data <= in_data_12_9;
			10'b0110001010 : out_data <= in_data_12_10;
			10'b0110001011 : out_data <= in_data_12_11;
			10'b0110001100 : out_data <= in_data_12_12;
			10'b0110001101 : out_data <= in_data_12_13;
			10'b0110001110 : out_data <= in_data_12_14;
			10'b0110001111 : out_data <= in_data_12_15;
			10'b0110010000 : out_data <= in_data_12_16;
			10'b0110010001 : out_data <= in_data_12_17;
			10'b0110010010 : out_data <= in_data_12_18;
			10'b0110010011 : out_data <= in_data_12_19;
			10'b0110010100 : out_data <= in_data_12_20;
			10'b0110010101 : out_data <= in_data_12_21;
			10'b0110010110 : out_data <= in_data_12_22;
			10'b0110010111 : out_data <= in_data_12_23;
			10'b0110011000 : out_data <= in_data_12_24;
			10'b0110011001 : out_data <= in_data_12_25;
			10'b0110011010 : out_data <= in_data_12_26;
			10'b0110011011 : out_data <= in_data_12_27;
			10'b0110011100 : out_data <= in_data_12_28;
			10'b0110011101 : out_data <= in_data_12_29;
			10'b0110011110 : out_data <= in_data_12_30;
			10'b0110011111 : out_data <= in_data_12_31;
			10'b0110100000 : out_data <= in_data_13_0;
			10'b0110100001 : out_data <= in_data_13_1;
			10'b0110100010 : out_data <= in_data_13_2;
			10'b0110100011 : out_data <= in_data_13_3;
			10'b0110100100 : out_data <= in_data_13_4;
			10'b0110100101 : out_data <= in_data_13_5;
			10'b0110100110 : out_data <= in_data_13_6;
			10'b0110100111 : out_data <= in_data_13_7;
			10'b0110101000 : out_data <= in_data_13_8;
			10'b0110101001 : out_data <= in_data_13_9;
			10'b0110101010 : out_data <= in_data_13_10;
			10'b0110101011 : out_data <= in_data_13_11;
			10'b0110101100 : out_data <= in_data_13_12;
			10'b0110101101 : out_data <= in_data_13_13;
			10'b0110101110 : out_data <= in_data_13_14;
			10'b0110101111 : out_data <= in_data_13_15;
			10'b0110110000 : out_data <= in_data_13_16;
			10'b0110110001 : out_data <= in_data_13_17;
			10'b0110110010 : out_data <= in_data_13_18;
			10'b0110110011 : out_data <= in_data_13_19;
			10'b0110110100 : out_data <= in_data_13_20;
			10'b0110110101 : out_data <= in_data_13_21;
			10'b0110110110 : out_data <= in_data_13_22;
			10'b0110110111 : out_data <= in_data_13_23;
			10'b0110111000 : out_data <= in_data_13_24;
			10'b0110111001 : out_data <= in_data_13_25;
			10'b0110111010 : out_data <= in_data_13_26;
			10'b0110111011 : out_data <= in_data_13_27;
			10'b0110111100 : out_data <= in_data_13_28;
			10'b0110111101 : out_data <= in_data_13_29;
			10'b0110111110 : out_data <= in_data_13_30;
			10'b0110111111 : out_data <= in_data_13_31;
			10'b0111000000 : out_data <= in_data_14_0;
			10'b0111000001 : out_data <= in_data_14_1;
			10'b0111000010 : out_data <= in_data_14_2;
			10'b0111000011 : out_data <= in_data_14_3;
			10'b0111000100 : out_data <= in_data_14_4;
			10'b0111000101 : out_data <= in_data_14_5;
			10'b0111000110 : out_data <= in_data_14_6;
			10'b0111000111 : out_data <= in_data_14_7;
			10'b0111001000 : out_data <= in_data_14_8;
			10'b0111001001 : out_data <= in_data_14_9;
			10'b0111001010 : out_data <= in_data_14_10;
			10'b0111001011 : out_data <= in_data_14_11;
			10'b0111001100 : out_data <= in_data_14_12;
			10'b0111001101 : out_data <= in_data_14_13;
			10'b0111001110 : out_data <= in_data_14_14;
			10'b0111001111 : out_data <= in_data_14_15;
			10'b0111010000 : out_data <= in_data_14_16;
			10'b0111010001 : out_data <= in_data_14_17;
			10'b0111010010 : out_data <= in_data_14_18;
			10'b0111010011 : out_data <= in_data_14_19;
			10'b0111010100 : out_data <= in_data_14_20;
			10'b0111010101 : out_data <= in_data_14_21;
			10'b0111010110 : out_data <= in_data_14_22;
			10'b0111010111 : out_data <= in_data_14_23;
			10'b0111011000 : out_data <= in_data_14_24;
			10'b0111011001 : out_data <= in_data_14_25;
			10'b0111011010 : out_data <= in_data_14_26;
			10'b0111011011 : out_data <= in_data_14_27;
			10'b0111011100 : out_data <= in_data_14_28;
			10'b0111011101 : out_data <= in_data_14_29;
			10'b0111011110 : out_data <= in_data_14_30;
			10'b0111011111 : out_data <= in_data_14_31;
			10'b0111100000 : out_data <= in_data_15_0;
			10'b0111100001 : out_data <= in_data_15_1;
			10'b0111100010 : out_data <= in_data_15_2;
			10'b0111100011 : out_data <= in_data_15_3;
			10'b0111100100 : out_data <= in_data_15_4;
			10'b0111100101 : out_data <= in_data_15_5;
			10'b0111100110 : out_data <= in_data_15_6;
			10'b0111100111 : out_data <= in_data_15_7;
			10'b0111101000 : out_data <= in_data_15_8;
			10'b0111101001 : out_data <= in_data_15_9;
			10'b0111101010 : out_data <= in_data_15_10;
			10'b0111101011 : out_data <= in_data_15_11;
			10'b0111101100 : out_data <= in_data_15_12;
			10'b0111101101 : out_data <= in_data_15_13;
			10'b0111101110 : out_data <= in_data_15_14;
			10'b0111101111 : out_data <= in_data_15_15;
			10'b0111110000 : out_data <= in_data_15_16;
			10'b0111110001 : out_data <= in_data_15_17;
			10'b0111110010 : out_data <= in_data_15_18;
			10'b0111110011 : out_data <= in_data_15_19;
			10'b0111110100 : out_data <= in_data_15_20;
			10'b0111110101 : out_data <= in_data_15_21;
			10'b0111110110 : out_data <= in_data_15_22;
			10'b0111110111 : out_data <= in_data_15_23;
			10'b0111111000 : out_data <= in_data_15_24;
			10'b0111111001 : out_data <= in_data_15_25;
			10'b0111111010 : out_data <= in_data_15_26;
			10'b0111111011 : out_data <= in_data_15_27;
			10'b0111111100 : out_data <= in_data_15_28;
			10'b0111111101 : out_data <= in_data_15_29;
			10'b0111111110 : out_data <= in_data_15_30;
			10'b0111111111 : out_data <= in_data_15_31;
			10'b1000000000 : out_data <= in_data_16_0;
			10'b1000000001 : out_data <= in_data_16_1;
			10'b1000000010 : out_data <= in_data_16_2;
			10'b1000000011 : out_data <= in_data_16_3;
			10'b1000000100 : out_data <= in_data_16_4;
			10'b1000000101 : out_data <= in_data_16_5;
			10'b1000000110 : out_data <= in_data_16_6;
			10'b1000000111 : out_data <= in_data_16_7;
			10'b1000001000 : out_data <= in_data_16_8;
			10'b1000001001 : out_data <= in_data_16_9;
			10'b1000001010 : out_data <= in_data_16_10;
			10'b1000001011 : out_data <= in_data_16_11;
			10'b1000001100 : out_data <= in_data_16_12;
			10'b1000001101 : out_data <= in_data_16_13;
			10'b1000001110 : out_data <= in_data_16_14;
			10'b1000001111 : out_data <= in_data_16_15;
			10'b1000010000 : out_data <= in_data_16_16;
			10'b1000010001 : out_data <= in_data_16_17;
			10'b1000010010 : out_data <= in_data_16_18;
			10'b1000010011 : out_data <= in_data_16_19;
			10'b1000010100 : out_data <= in_data_16_20;
			10'b1000010101 : out_data <= in_data_16_21;
			10'b1000010110 : out_data <= in_data_16_22;
			10'b1000010111 : out_data <= in_data_16_23;
			10'b1000011000 : out_data <= in_data_16_24;
			10'b1000011001 : out_data <= in_data_16_25;
			10'b1000011010 : out_data <= in_data_16_26;
			10'b1000011011 : out_data <= in_data_16_27;
			10'b1000011100 : out_data <= in_data_16_28;
			10'b1000011101 : out_data <= in_data_16_29;
			10'b1000011110 : out_data <= in_data_16_30;
			10'b1000011111 : out_data <= in_data_16_31;
			10'b1000100000 : out_data <= in_data_17_0;
			10'b1000100001 : out_data <= in_data_17_1;
			10'b1000100010 : out_data <= in_data_17_2;
			10'b1000100011 : out_data <= in_data_17_3;
			10'b1000100100 : out_data <= in_data_17_4;
			10'b1000100101 : out_data <= in_data_17_5;
			10'b1000100110 : out_data <= in_data_17_6;
			10'b1000100111 : out_data <= in_data_17_7;
			10'b1000101000 : out_data <= in_data_17_8;
			10'b1000101001 : out_data <= in_data_17_9;
			10'b1000101010 : out_data <= in_data_17_10;
			10'b1000101011 : out_data <= in_data_17_11;
			10'b1000101100 : out_data <= in_data_17_12;
			10'b1000101101 : out_data <= in_data_17_13;
			10'b1000101110 : out_data <= in_data_17_14;
			10'b1000101111 : out_data <= in_data_17_15;
			10'b1000110000 : out_data <= in_data_17_16;
			10'b1000110001 : out_data <= in_data_17_17;
			10'b1000110010 : out_data <= in_data_17_18;
			10'b1000110011 : out_data <= in_data_17_19;
			10'b1000110100 : out_data <= in_data_17_20;
			10'b1000110101 : out_data <= in_data_17_21;
			10'b1000110110 : out_data <= in_data_17_22;
			10'b1000110111 : out_data <= in_data_17_23;
			10'b1000111000 : out_data <= in_data_17_24;
			10'b1000111001 : out_data <= in_data_17_25;
			10'b1000111010 : out_data <= in_data_17_26;
			10'b1000111011 : out_data <= in_data_17_27;
			10'b1000111100 : out_data <= in_data_17_28;
			10'b1000111101 : out_data <= in_data_17_29;
			10'b1000111110 : out_data <= in_data_17_30;
			10'b1000111111 : out_data <= in_data_17_31;
			10'b1001000000 : out_data <= in_data_18_0;
			10'b1001000001 : out_data <= in_data_18_1;
			10'b1001000010 : out_data <= in_data_18_2;
			10'b1001000011 : out_data <= in_data_18_3;
			10'b1001000100 : out_data <= in_data_18_4;
			10'b1001000101 : out_data <= in_data_18_5;
			10'b1001000110 : out_data <= in_data_18_6;
			10'b1001000111 : out_data <= in_data_18_7;
			10'b1001001000 : out_data <= in_data_18_8;
			10'b1001001001 : out_data <= in_data_18_9;
			10'b1001001010 : out_data <= in_data_18_10;
			10'b1001001011 : out_data <= in_data_18_11;
			10'b1001001100 : out_data <= in_data_18_12;
			10'b1001001101 : out_data <= in_data_18_13;
			10'b1001001110 : out_data <= in_data_18_14;
			10'b1001001111 : out_data <= in_data_18_15;
			10'b1001010000 : out_data <= in_data_18_16;
			10'b1001010001 : out_data <= in_data_18_17;
			10'b1001010010 : out_data <= in_data_18_18;
			10'b1001010011 : out_data <= in_data_18_19;
			10'b1001010100 : out_data <= in_data_18_20;
			10'b1001010101 : out_data <= in_data_18_21;
			10'b1001010110 : out_data <= in_data_18_22;
			10'b1001010111 : out_data <= in_data_18_23;
			10'b1001011000 : out_data <= in_data_18_24;
			10'b1001011001 : out_data <= in_data_18_25;
			10'b1001011010 : out_data <= in_data_18_26;
			10'b1001011011 : out_data <= in_data_18_27;
			10'b1001011100 : out_data <= in_data_18_28;
			10'b1001011101 : out_data <= in_data_18_29;
			10'b1001011110 : out_data <= in_data_18_30;
			10'b1001011111 : out_data <= in_data_18_31;
			10'b1001100000 : out_data <= in_data_19_0;
			10'b1001100001 : out_data <= in_data_19_1;
			10'b1001100010 : out_data <= in_data_19_2;
			10'b1001100011 : out_data <= in_data_19_3;
			10'b1001100100 : out_data <= in_data_19_4;
			10'b1001100101 : out_data <= in_data_19_5;
			10'b1001100110 : out_data <= in_data_19_6;
			10'b1001100111 : out_data <= in_data_19_7;
			10'b1001101000 : out_data <= in_data_19_8;
			10'b1001101001 : out_data <= in_data_19_9;
			10'b1001101010 : out_data <= in_data_19_10;
			10'b1001101011 : out_data <= in_data_19_11;
			10'b1001101100 : out_data <= in_data_19_12;
			10'b1001101101 : out_data <= in_data_19_13;
			10'b1001101110 : out_data <= in_data_19_14;
			10'b1001101111 : out_data <= in_data_19_15;
			10'b1001110000 : out_data <= in_data_19_16;
			10'b1001110001 : out_data <= in_data_19_17;
			10'b1001110010 : out_data <= in_data_19_18;
			10'b1001110011 : out_data <= in_data_19_19;
			10'b1001110100 : out_data <= in_data_19_20;
			10'b1001110101 : out_data <= in_data_19_21;
			10'b1001110110 : out_data <= in_data_19_22;
			10'b1001110111 : out_data <= in_data_19_23;
			10'b1001111000 : out_data <= in_data_19_24;
			10'b1001111001 : out_data <= in_data_19_25;
			10'b1001111010 : out_data <= in_data_19_26;
			10'b1001111011 : out_data <= in_data_19_27;
			10'b1001111100 : out_data <= in_data_19_28;
			10'b1001111101 : out_data <= in_data_19_29;
			10'b1001111110 : out_data <= in_data_19_30;
			10'b1001111111 : out_data <= in_data_19_31;
			10'b1010000000 : out_data <= in_data_20_0;
			10'b1010000001 : out_data <= in_data_20_1;
			10'b1010000010 : out_data <= in_data_20_2;
			10'b1010000011 : out_data <= in_data_20_3;
			10'b1010000100 : out_data <= in_data_20_4;
			10'b1010000101 : out_data <= in_data_20_5;
			10'b1010000110 : out_data <= in_data_20_6;
			10'b1010000111 : out_data <= in_data_20_7;
			10'b1010001000 : out_data <= in_data_20_8;
			10'b1010001001 : out_data <= in_data_20_9;
			10'b1010001010 : out_data <= in_data_20_10;
			10'b1010001011 : out_data <= in_data_20_11;
			10'b1010001100 : out_data <= in_data_20_12;
			10'b1010001101 : out_data <= in_data_20_13;
			10'b1010001110 : out_data <= in_data_20_14;
			10'b1010001111 : out_data <= in_data_20_15;
			10'b1010010000 : out_data <= in_data_20_16;
			10'b1010010001 : out_data <= in_data_20_17;
			10'b1010010010 : out_data <= in_data_20_18;
			10'b1010010011 : out_data <= in_data_20_19;
			10'b1010010100 : out_data <= in_data_20_20;
			10'b1010010101 : out_data <= in_data_20_21;
			10'b1010010110 : out_data <= in_data_20_22;
			10'b1010010111 : out_data <= in_data_20_23;
			10'b1010011000 : out_data <= in_data_20_24;
			10'b1010011001 : out_data <= in_data_20_25;
			10'b1010011010 : out_data <= in_data_20_26;
			10'b1010011011 : out_data <= in_data_20_27;
			10'b1010011100 : out_data <= in_data_20_28;
			10'b1010011101 : out_data <= in_data_20_29;
			10'b1010011110 : out_data <= in_data_20_30;
			10'b1010011111 : out_data <= in_data_20_31;
			10'b1010100000 : out_data <= in_data_21_0;
			10'b1010100001 : out_data <= in_data_21_1;
			10'b1010100010 : out_data <= in_data_21_2;
			10'b1010100011 : out_data <= in_data_21_3;
			10'b1010100100 : out_data <= in_data_21_4;
			10'b1010100101 : out_data <= in_data_21_5;
			10'b1010100110 : out_data <= in_data_21_6;
			10'b1010100111 : out_data <= in_data_21_7;
			10'b1010101000 : out_data <= in_data_21_8;
			10'b1010101001 : out_data <= in_data_21_9;
			10'b1010101010 : out_data <= in_data_21_10;
			10'b1010101011 : out_data <= in_data_21_11;
			10'b1010101100 : out_data <= in_data_21_12;
			10'b1010101101 : out_data <= in_data_21_13;
			10'b1010101110 : out_data <= in_data_21_14;
			10'b1010101111 : out_data <= in_data_21_15;
			10'b1010110000 : out_data <= in_data_21_16;
			10'b1010110001 : out_data <= in_data_21_17;
			10'b1010110010 : out_data <= in_data_21_18;
			10'b1010110011 : out_data <= in_data_21_19;
			10'b1010110100 : out_data <= in_data_21_20;
			10'b1010110101 : out_data <= in_data_21_21;
			10'b1010110110 : out_data <= in_data_21_22;
			10'b1010110111 : out_data <= in_data_21_23;
			10'b1010111000 : out_data <= in_data_21_24;
			10'b1010111001 : out_data <= in_data_21_25;
			10'b1010111010 : out_data <= in_data_21_26;
			10'b1010111011 : out_data <= in_data_21_27;
			10'b1010111100 : out_data <= in_data_21_28;
			10'b1010111101 : out_data <= in_data_21_29;
			10'b1010111110 : out_data <= in_data_21_30;
			10'b1010111111 : out_data <= in_data_21_31;
			10'b1011000000 : out_data <= in_data_22_0;
			10'b1011000001 : out_data <= in_data_22_1;
			10'b1011000010 : out_data <= in_data_22_2;
			10'b1011000011 : out_data <= in_data_22_3;
			10'b1011000100 : out_data <= in_data_22_4;
			10'b1011000101 : out_data <= in_data_22_5;
			10'b1011000110 : out_data <= in_data_22_6;
			10'b1011000111 : out_data <= in_data_22_7;
			10'b1011001000 : out_data <= in_data_22_8;
			10'b1011001001 : out_data <= in_data_22_9;
			10'b1011001010 : out_data <= in_data_22_10;
			10'b1011001011 : out_data <= in_data_22_11;
			10'b1011001100 : out_data <= in_data_22_12;
			10'b1011001101 : out_data <= in_data_22_13;
			10'b1011001110 : out_data <= in_data_22_14;
			10'b1011001111 : out_data <= in_data_22_15;
			10'b1011010000 : out_data <= in_data_22_16;
			10'b1011010001 : out_data <= in_data_22_17;
			10'b1011010010 : out_data <= in_data_22_18;
			10'b1011010011 : out_data <= in_data_22_19;
			10'b1011010100 : out_data <= in_data_22_20;
			10'b1011010101 : out_data <= in_data_22_21;
			10'b1011010110 : out_data <= in_data_22_22;
			10'b1011010111 : out_data <= in_data_22_23;
			10'b1011011000 : out_data <= in_data_22_24;
			10'b1011011001 : out_data <= in_data_22_25;
			10'b1011011010 : out_data <= in_data_22_26;
			10'b1011011011 : out_data <= in_data_22_27;
			10'b1011011100 : out_data <= in_data_22_28;
			10'b1011011101 : out_data <= in_data_22_29;
			10'b1011011110 : out_data <= in_data_22_30;
			10'b1011011111 : out_data <= in_data_22_31;
			10'b1011100000 : out_data <= in_data_23_0;
			10'b1011100001 : out_data <= in_data_23_1;
			10'b1011100010 : out_data <= in_data_23_2;
			10'b1011100011 : out_data <= in_data_23_3;
			10'b1011100100 : out_data <= in_data_23_4;
			10'b1011100101 : out_data <= in_data_23_5;
			10'b1011100110 : out_data <= in_data_23_6;
			10'b1011100111 : out_data <= in_data_23_7;
			10'b1011101000 : out_data <= in_data_23_8;
			10'b1011101001 : out_data <= in_data_23_9;
			10'b1011101010 : out_data <= in_data_23_10;
			10'b1011101011 : out_data <= in_data_23_11;
			10'b1011101100 : out_data <= in_data_23_12;
			10'b1011101101 : out_data <= in_data_23_13;
			10'b1011101110 : out_data <= in_data_23_14;
			10'b1011101111 : out_data <= in_data_23_15;
			10'b1011110000 : out_data <= in_data_23_16;
			10'b1011110001 : out_data <= in_data_23_17;
			10'b1011110010 : out_data <= in_data_23_18;
			10'b1011110011 : out_data <= in_data_23_19;
			10'b1011110100 : out_data <= in_data_23_20;
			10'b1011110101 : out_data <= in_data_23_21;
			10'b1011110110 : out_data <= in_data_23_22;
			10'b1011110111 : out_data <= in_data_23_23;
			10'b1011111000 : out_data <= in_data_23_24;
			10'b1011111001 : out_data <= in_data_23_25;
			10'b1011111010 : out_data <= in_data_23_26;
			10'b1011111011 : out_data <= in_data_23_27;
			10'b1011111100 : out_data <= in_data_23_28;
			10'b1011111101 : out_data <= in_data_23_29;
			10'b1011111110 : out_data <= in_data_23_30;
			10'b1011111111 : out_data <= in_data_23_31;
			10'b1100000000 : out_data <= in_data_24_0;
			10'b1100000001 : out_data <= in_data_24_1;
			10'b1100000010 : out_data <= in_data_24_2;
			10'b1100000011 : out_data <= in_data_24_3;
			10'b1100000100 : out_data <= in_data_24_4;
			10'b1100000101 : out_data <= in_data_24_5;
			10'b1100000110 : out_data <= in_data_24_6;
			10'b1100000111 : out_data <= in_data_24_7;
			10'b1100001000 : out_data <= in_data_24_8;
			10'b1100001001 : out_data <= in_data_24_9;
			10'b1100001010 : out_data <= in_data_24_10;
			10'b1100001011 : out_data <= in_data_24_11;
			10'b1100001100 : out_data <= in_data_24_12;
			10'b1100001101 : out_data <= in_data_24_13;
			10'b1100001110 : out_data <= in_data_24_14;
			10'b1100001111 : out_data <= in_data_24_15;
			10'b1100010000 : out_data <= in_data_24_16;
			10'b1100010001 : out_data <= in_data_24_17;
			10'b1100010010 : out_data <= in_data_24_18;
			10'b1100010011 : out_data <= in_data_24_19;
			10'b1100010100 : out_data <= in_data_24_20;
			10'b1100010101 : out_data <= in_data_24_21;
			10'b1100010110 : out_data <= in_data_24_22;
			10'b1100010111 : out_data <= in_data_24_23;
			10'b1100011000 : out_data <= in_data_24_24;
			10'b1100011001 : out_data <= in_data_24_25;
			10'b1100011010 : out_data <= in_data_24_26;
			10'b1100011011 : out_data <= in_data_24_27;
			10'b1100011100 : out_data <= in_data_24_28;
			10'b1100011101 : out_data <= in_data_24_29;
			10'b1100011110 : out_data <= in_data_24_30;
			10'b1100011111 : out_data <= in_data_24_31;
			10'b1100100000 : out_data <= in_data_25_0;
			10'b1100100001 : out_data <= in_data_25_1;
			10'b1100100010 : out_data <= in_data_25_2;
			10'b1100100011 : out_data <= in_data_25_3;
			10'b1100100100 : out_data <= in_data_25_4;
			10'b1100100101 : out_data <= in_data_25_5;
			10'b1100100110 : out_data <= in_data_25_6;
			10'b1100100111 : out_data <= in_data_25_7;
			10'b1100101000 : out_data <= in_data_25_8;
			10'b1100101001 : out_data <= in_data_25_9;
			10'b1100101010 : out_data <= in_data_25_10;
			10'b1100101011 : out_data <= in_data_25_11;
			10'b1100101100 : out_data <= in_data_25_12;
			10'b1100101101 : out_data <= in_data_25_13;
			10'b1100101110 : out_data <= in_data_25_14;
			10'b1100101111 : out_data <= in_data_25_15;
			10'b1100110000 : out_data <= in_data_25_16;
			10'b1100110001 : out_data <= in_data_25_17;
			10'b1100110010 : out_data <= in_data_25_18;
			10'b1100110011 : out_data <= in_data_25_19;
			10'b1100110100 : out_data <= in_data_25_20;
			10'b1100110101 : out_data <= in_data_25_21;
			10'b1100110110 : out_data <= in_data_25_22;
			10'b1100110111 : out_data <= in_data_25_23;
			10'b1100111000 : out_data <= in_data_25_24;
			10'b1100111001 : out_data <= in_data_25_25;
			10'b1100111010 : out_data <= in_data_25_26;
			10'b1100111011 : out_data <= in_data_25_27;
			10'b1100111100 : out_data <= in_data_25_28;
			10'b1100111101 : out_data <= in_data_25_29;
			10'b1100111110 : out_data <= in_data_25_30;
			10'b1100111111 : out_data <= in_data_25_31;
			10'b1101000000 : out_data <= in_data_26_0;
			10'b1101000001 : out_data <= in_data_26_1;
			10'b1101000010 : out_data <= in_data_26_2;
			10'b1101000011 : out_data <= in_data_26_3;
			10'b1101000100 : out_data <= in_data_26_4;
			10'b1101000101 : out_data <= in_data_26_5;
			10'b1101000110 : out_data <= in_data_26_6;
			10'b1101000111 : out_data <= in_data_26_7;
			10'b1101001000 : out_data <= in_data_26_8;
			10'b1101001001 : out_data <= in_data_26_9;
			10'b1101001010 : out_data <= in_data_26_10;
			10'b1101001011 : out_data <= in_data_26_11;
			10'b1101001100 : out_data <= in_data_26_12;
			10'b1101001101 : out_data <= in_data_26_13;
			10'b1101001110 : out_data <= in_data_26_14;
			10'b1101001111 : out_data <= in_data_26_15;
			10'b1101010000 : out_data <= in_data_26_16;
			10'b1101010001 : out_data <= in_data_26_17;
			10'b1101010010 : out_data <= in_data_26_18;
			10'b1101010011 : out_data <= in_data_26_19;
			10'b1101010100 : out_data <= in_data_26_20;
			10'b1101010101 : out_data <= in_data_26_21;
			10'b1101010110 : out_data <= in_data_26_22;
			10'b1101010111 : out_data <= in_data_26_23;
			10'b1101011000 : out_data <= in_data_26_24;
			10'b1101011001 : out_data <= in_data_26_25;
			10'b1101011010 : out_data <= in_data_26_26;
			10'b1101011011 : out_data <= in_data_26_27;
			10'b1101011100 : out_data <= in_data_26_28;
			10'b1101011101 : out_data <= in_data_26_29;
			10'b1101011110 : out_data <= in_data_26_30;
			10'b1101011111 : out_data <= in_data_26_31;
			10'b1101100000 : out_data <= in_data_27_0;
			10'b1101100001 : out_data <= in_data_27_1;
			10'b1101100010 : out_data <= in_data_27_2;
			10'b1101100011 : out_data <= in_data_27_3;
			10'b1101100100 : out_data <= in_data_27_4;
			10'b1101100101 : out_data <= in_data_27_5;
			10'b1101100110 : out_data <= in_data_27_6;
			10'b1101100111 : out_data <= in_data_27_7;
			10'b1101101000 : out_data <= in_data_27_8;
			10'b1101101001 : out_data <= in_data_27_9;
			10'b1101101010 : out_data <= in_data_27_10;
			10'b1101101011 : out_data <= in_data_27_11;
			10'b1101101100 : out_data <= in_data_27_12;
			10'b1101101101 : out_data <= in_data_27_13;
			10'b1101101110 : out_data <= in_data_27_14;
			10'b1101101111 : out_data <= in_data_27_15;
			10'b1101110000 : out_data <= in_data_27_16;
			10'b1101110001 : out_data <= in_data_27_17;
			10'b1101110010 : out_data <= in_data_27_18;
			10'b1101110011 : out_data <= in_data_27_19;
			10'b1101110100 : out_data <= in_data_27_20;
			10'b1101110101 : out_data <= in_data_27_21;
			10'b1101110110 : out_data <= in_data_27_22;
			10'b1101110111 : out_data <= in_data_27_23;
			10'b1101111000 : out_data <= in_data_27_24;
			10'b1101111001 : out_data <= in_data_27_25;
			10'b1101111010 : out_data <= in_data_27_26;
			10'b1101111011 : out_data <= in_data_27_27;
			10'b1101111100 : out_data <= in_data_27_28;
			10'b1101111101 : out_data <= in_data_27_29;
			10'b1101111110 : out_data <= in_data_27_30;
			10'b1101111111 : out_data <= in_data_27_31;
			10'b1110000000 : out_data <= in_data_28_0;
			10'b1110000001 : out_data <= in_data_28_1;
			10'b1110000010 : out_data <= in_data_28_2;
			10'b1110000011 : out_data <= in_data_28_3;
			10'b1110000100 : out_data <= in_data_28_4;
			10'b1110000101 : out_data <= in_data_28_5;
			10'b1110000110 : out_data <= in_data_28_6;
			10'b1110000111 : out_data <= in_data_28_7;
			10'b1110001000 : out_data <= in_data_28_8;
			10'b1110001001 : out_data <= in_data_28_9;
			10'b1110001010 : out_data <= in_data_28_10;
			10'b1110001011 : out_data <= in_data_28_11;
			10'b1110001100 : out_data <= in_data_28_12;
			10'b1110001101 : out_data <= in_data_28_13;
			10'b1110001110 : out_data <= in_data_28_14;
			10'b1110001111 : out_data <= in_data_28_15;
			10'b1110010000 : out_data <= in_data_28_16;
			10'b1110010001 : out_data <= in_data_28_17;
			10'b1110010010 : out_data <= in_data_28_18;
			10'b1110010011 : out_data <= in_data_28_19;
			10'b1110010100 : out_data <= in_data_28_20;
			10'b1110010101 : out_data <= in_data_28_21;
			10'b1110010110 : out_data <= in_data_28_22;
			10'b1110010111 : out_data <= in_data_28_23;
			10'b1110011000 : out_data <= in_data_28_24;
			10'b1110011001 : out_data <= in_data_28_25;
			10'b1110011010 : out_data <= in_data_28_26;
			10'b1110011011 : out_data <= in_data_28_27;
			10'b1110011100 : out_data <= in_data_28_28;
			10'b1110011101 : out_data <= in_data_28_29;
			10'b1110011110 : out_data <= in_data_28_30;
			10'b1110011111 : out_data <= in_data_28_31;
			10'b1110100000 : out_data <= in_data_29_0;
			10'b1110100001 : out_data <= in_data_29_1;
			10'b1110100010 : out_data <= in_data_29_2;
			10'b1110100011 : out_data <= in_data_29_3;
			10'b1110100100 : out_data <= in_data_29_4;
			10'b1110100101 : out_data <= in_data_29_5;
			10'b1110100110 : out_data <= in_data_29_6;
			10'b1110100111 : out_data <= in_data_29_7;
			10'b1110101000 : out_data <= in_data_29_8;
			10'b1110101001 : out_data <= in_data_29_9;
			10'b1110101010 : out_data <= in_data_29_10;
			10'b1110101011 : out_data <= in_data_29_11;
			10'b1110101100 : out_data <= in_data_29_12;
			10'b1110101101 : out_data <= in_data_29_13;
			10'b1110101110 : out_data <= in_data_29_14;
			10'b1110101111 : out_data <= in_data_29_15;
			10'b1110110000 : out_data <= in_data_29_16;
			10'b1110110001 : out_data <= in_data_29_17;
			10'b1110110010 : out_data <= in_data_29_18;
			10'b1110110011 : out_data <= in_data_29_19;
			10'b1110110100 : out_data <= in_data_29_20;
			10'b1110110101 : out_data <= in_data_29_21;
			10'b1110110110 : out_data <= in_data_29_22;
			10'b1110110111 : out_data <= in_data_29_23;
			10'b1110111000 : out_data <= in_data_29_24;
			10'b1110111001 : out_data <= in_data_29_25;
			10'b1110111010 : out_data <= in_data_29_26;
			10'b1110111011 : out_data <= in_data_29_27;
			10'b1110111100 : out_data <= in_data_29_28;
			10'b1110111101 : out_data <= in_data_29_29;
			10'b1110111110 : out_data <= in_data_29_30;
			10'b1110111111 : out_data <= in_data_29_31;
			10'b1111000000 : out_data <= in_data_30_0;
			10'b1111000001 : out_data <= in_data_30_1;
			10'b1111000010 : out_data <= in_data_30_2;
			10'b1111000011 : out_data <= in_data_30_3;
			10'b1111000100 : out_data <= in_data_30_4;
			10'b1111000101 : out_data <= in_data_30_5;
			10'b1111000110 : out_data <= in_data_30_6;
			10'b1111000111 : out_data <= in_data_30_7;
			10'b1111001000 : out_data <= in_data_30_8;
			10'b1111001001 : out_data <= in_data_30_9;
			10'b1111001010 : out_data <= in_data_30_10;
			10'b1111001011 : out_data <= in_data_30_11;
			10'b1111001100 : out_data <= in_data_30_12;
			10'b1111001101 : out_data <= in_data_30_13;
			10'b1111001110 : out_data <= in_data_30_14;
			10'b1111001111 : out_data <= in_data_30_15;
			10'b1111010000 : out_data <= in_data_30_16;
			10'b1111010001 : out_data <= in_data_30_17;
			10'b1111010010 : out_data <= in_data_30_18;
			10'b1111010011 : out_data <= in_data_30_19;
			10'b1111010100 : out_data <= in_data_30_20;
			10'b1111010101 : out_data <= in_data_30_21;
			10'b1111010110 : out_data <= in_data_30_22;
			10'b1111010111 : out_data <= in_data_30_23;
			10'b1111011000 : out_data <= in_data_30_24;
			10'b1111011001 : out_data <= in_data_30_25;
			10'b1111011010 : out_data <= in_data_30_26;
			10'b1111011011 : out_data <= in_data_30_27;
			10'b1111011100 : out_data <= in_data_30_28;
			10'b1111011101 : out_data <= in_data_30_29;
			10'b1111011110 : out_data <= in_data_30_30;
			10'b1111011111 : out_data <= in_data_30_31;
			10'b1111100000 : out_data <= in_data_31_0;
			10'b1111100001 : out_data <= in_data_31_1;
			10'b1111100010 : out_data <= in_data_31_2;
			10'b1111100011 : out_data <= in_data_31_3;
			10'b1111100100 : out_data <= in_data_31_4;
			10'b1111100101 : out_data <= in_data_31_5;
			10'b1111100110 : out_data <= in_data_31_6;
			10'b1111100111 : out_data <= in_data_31_7;
			10'b1111101000 : out_data <= in_data_31_8;
			10'b1111101001 : out_data <= in_data_31_9;
			10'b1111101010 : out_data <= in_data_31_10;
			10'b1111101011 : out_data <= in_data_31_11;
			10'b1111101100 : out_data <= in_data_31_12;
			10'b1111101101 : out_data <= in_data_31_13;
			10'b1111101110 : out_data <= in_data_31_14;
			10'b1111101111 : out_data <= in_data_31_15;
			10'b1111110000 : out_data <= in_data_31_16;
			10'b1111110001 : out_data <= in_data_31_17;
			10'b1111110010 : out_data <= in_data_31_18;
			10'b1111110011 : out_data <= in_data_31_19;
			10'b1111110100 : out_data <= in_data_31_20;
			10'b1111110101 : out_data <= in_data_31_21;
			10'b1111110110 : out_data <= in_data_31_22;
			10'b1111110111 : out_data <= in_data_31_23;
			10'b1111111000 : out_data <= in_data_31_24;
			10'b1111111001 : out_data <= in_data_31_25;
			10'b1111111010 : out_data <= in_data_31_26;
			10'b1111111011 : out_data <= in_data_31_27;
			10'b1111111100 : out_data <= in_data_31_28;
			10'b1111111101 : out_data <= in_data_31_29;
			10'b1111111110 : out_data <= in_data_31_30;
			10'b1111111111 : out_data <= in_data_31_31;
  endcase
end

endmodule
