`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: TODO
// Engineer: TODO
//
// Create Date: 2024-09-06 17:06:52.512677
// Target Devices: TODO
// Tool Versions: TODO
// Description: TODO
//
// Additional Comments:
////////////////////////////////////////////////////////////////////////////////
module systolic_array_32x32 #(parameter DEPTH=8, DATA_WIDTH=16, OUT_SELECT_WIDTH=10) (
	input clk, rstn,
	input r_en, w_en,
	input [4:0] row_select,
	input [4:0] col_select,
	input [OUT_SELECT_WIDTH-1:0] out_select,
	input signed [DATA_WIDTH-1:0] in_row,
	input signed [DATA_WIDTH-1:0] in_col,
	output signed [DATA_WIDTH-1:0] mux_data_out,
	output row_fifo_0_full,
	output row_fifo_0_empty,
	output row_fifo_1_full,
	output row_fifo_1_empty,
	output row_fifo_2_full,
	output row_fifo_2_empty,
	output row_fifo_3_full,
	output row_fifo_3_empty,
	output row_fifo_4_full,
	output row_fifo_4_empty,
	output row_fifo_5_full,
	output row_fifo_5_empty,
	output row_fifo_6_full,
	output row_fifo_6_empty,
	output row_fifo_7_full,
	output row_fifo_7_empty,
	output row_fifo_8_full,
	output row_fifo_8_empty,
	output row_fifo_9_full,
	output row_fifo_9_empty,
	output row_fifo_10_full,
	output row_fifo_10_empty,
	output row_fifo_11_full,
	output row_fifo_11_empty,
	output row_fifo_12_full,
	output row_fifo_12_empty,
	output row_fifo_13_full,
	output row_fifo_13_empty,
	output row_fifo_14_full,
	output row_fifo_14_empty,
	output row_fifo_15_full,
	output row_fifo_15_empty,
	output row_fifo_16_full,
	output row_fifo_16_empty,
	output row_fifo_17_full,
	output row_fifo_17_empty,
	output row_fifo_18_full,
	output row_fifo_18_empty,
	output row_fifo_19_full,
	output row_fifo_19_empty,
	output row_fifo_20_full,
	output row_fifo_20_empty,
	output row_fifo_21_full,
	output row_fifo_21_empty,
	output row_fifo_22_full,
	output row_fifo_22_empty,
	output row_fifo_23_full,
	output row_fifo_23_empty,
	output row_fifo_24_full,
	output row_fifo_24_empty,
	output row_fifo_25_full,
	output row_fifo_25_empty,
	output row_fifo_26_full,
	output row_fifo_26_empty,
	output row_fifo_27_full,
	output row_fifo_27_empty,
	output row_fifo_28_full,
	output row_fifo_28_empty,
	output row_fifo_29_full,
	output row_fifo_29_empty,
	output row_fifo_30_full,
	output row_fifo_30_empty,
	output row_fifo_31_full,
	output row_fifo_31_empty,
	output col_fifo_0_full,
	output col_fifo_0_empty,
	output col_fifo_1_full,
	output col_fifo_1_empty,
	output col_fifo_2_full,
	output col_fifo_2_empty,
	output col_fifo_3_full,
	output col_fifo_3_empty,
	output col_fifo_4_full,
	output col_fifo_4_empty,
	output col_fifo_5_full,
	output col_fifo_5_empty,
	output col_fifo_6_full,
	output col_fifo_6_empty,
	output col_fifo_7_full,
	output col_fifo_7_empty,
	output col_fifo_8_full,
	output col_fifo_8_empty,
	output col_fifo_9_full,
	output col_fifo_9_empty,
	output col_fifo_10_full,
	output col_fifo_10_empty,
	output col_fifo_11_full,
	output col_fifo_11_empty,
	output col_fifo_12_full,
	output col_fifo_12_empty,
	output col_fifo_13_full,
	output col_fifo_13_empty,
	output col_fifo_14_full,
	output col_fifo_14_empty,
	output col_fifo_15_full,
	output col_fifo_15_empty,
	output col_fifo_16_full,
	output col_fifo_16_empty,
	output col_fifo_17_full,
	output col_fifo_17_empty,
	output col_fifo_18_full,
	output col_fifo_18_empty,
	output col_fifo_19_full,
	output col_fifo_19_empty,
	output col_fifo_20_full,
	output col_fifo_20_empty,
	output col_fifo_21_full,
	output col_fifo_21_empty,
	output col_fifo_22_full,
	output col_fifo_22_empty,
	output col_fifo_23_full,
	output col_fifo_23_empty,
	output col_fifo_24_full,
	output col_fifo_24_empty,
	output col_fifo_25_full,
	output col_fifo_25_empty,
	output col_fifo_26_full,
	output col_fifo_26_empty,
	output col_fifo_27_full,
	output col_fifo_27_empty,
	output col_fifo_28_full,
	output col_fifo_28_empty,
	output col_fifo_29_full,
	output col_fifo_29_empty,
	output col_fifo_30_full,
	output col_fifo_30_empty,
	output col_fifo_31_full,
	output col_fifo_31_empty
);
	wire [DATA_WIDTH-1:0] row_demux_out_data_0;
	wire [DATA_WIDTH-1:0] row_demux_out_data_1;
	wire [DATA_WIDTH-1:0] row_demux_out_data_2;
	wire [DATA_WIDTH-1:0] row_demux_out_data_3;
	wire [DATA_WIDTH-1:0] row_demux_out_data_4;
	wire [DATA_WIDTH-1:0] row_demux_out_data_5;
	wire [DATA_WIDTH-1:0] row_demux_out_data_6;
	wire [DATA_WIDTH-1:0] row_demux_out_data_7;
	wire [DATA_WIDTH-1:0] row_demux_out_data_8;
	wire [DATA_WIDTH-1:0] row_demux_out_data_9;
	wire [DATA_WIDTH-1:0] row_demux_out_data_10;
	wire [DATA_WIDTH-1:0] row_demux_out_data_11;
	wire [DATA_WIDTH-1:0] row_demux_out_data_12;
	wire [DATA_WIDTH-1:0] row_demux_out_data_13;
	wire [DATA_WIDTH-1:0] row_demux_out_data_14;
	wire [DATA_WIDTH-1:0] row_demux_out_data_15;
	wire [DATA_WIDTH-1:0] row_demux_out_data_16;
	wire [DATA_WIDTH-1:0] row_demux_out_data_17;
	wire [DATA_WIDTH-1:0] row_demux_out_data_18;
	wire [DATA_WIDTH-1:0] row_demux_out_data_19;
	wire [DATA_WIDTH-1:0] row_demux_out_data_20;
	wire [DATA_WIDTH-1:0] row_demux_out_data_21;
	wire [DATA_WIDTH-1:0] row_demux_out_data_22;
	wire [DATA_WIDTH-1:0] row_demux_out_data_23;
	wire [DATA_WIDTH-1:0] row_demux_out_data_24;
	wire [DATA_WIDTH-1:0] row_demux_out_data_25;
	wire [DATA_WIDTH-1:0] row_demux_out_data_26;
	wire [DATA_WIDTH-1:0] row_demux_out_data_27;
	wire [DATA_WIDTH-1:0] row_demux_out_data_28;
	wire [DATA_WIDTH-1:0] row_demux_out_data_29;
	wire [DATA_WIDTH-1:0] row_demux_out_data_30;
	wire [DATA_WIDTH-1:0] row_demux_out_data_31;
	demux_1_to_32  row_demux (
		.select (row_select),
		.in_data (in_row),
		.out_data_0 (row_demux_out_data_0),
		.out_data_1 (row_demux_out_data_1),
		.out_data_2 (row_demux_out_data_2),
		.out_data_3 (row_demux_out_data_3),
		.out_data_4 (row_demux_out_data_4),
		.out_data_5 (row_demux_out_data_5),
		.out_data_6 (row_demux_out_data_6),
		.out_data_7 (row_demux_out_data_7),
		.out_data_8 (row_demux_out_data_8),
		.out_data_9 (row_demux_out_data_9),
		.out_data_10 (row_demux_out_data_10),
		.out_data_11 (row_demux_out_data_11),
		.out_data_12 (row_demux_out_data_12),
		.out_data_13 (row_demux_out_data_13),
		.out_data_14 (row_demux_out_data_14),
		.out_data_15 (row_demux_out_data_15),
		.out_data_16 (row_demux_out_data_16),
		.out_data_17 (row_demux_out_data_17),
		.out_data_18 (row_demux_out_data_18),
		.out_data_19 (row_demux_out_data_19),
		.out_data_20 (row_demux_out_data_20),
		.out_data_21 (row_demux_out_data_21),
		.out_data_22 (row_demux_out_data_22),
		.out_data_23 (row_demux_out_data_23),
		.out_data_24 (row_demux_out_data_24),
		.out_data_25 (row_demux_out_data_25),
		.out_data_26 (row_demux_out_data_26),
		.out_data_27 (row_demux_out_data_27),
		.out_data_28 (row_demux_out_data_28),
		.out_data_29 (row_demux_out_data_29),
		.out_data_30 (row_demux_out_data_30),
		.out_data_31 (row_demux_out_data_31)
	);
	wire [DATA_WIDTH-1:0] col_demux_out_data_0;
	wire [DATA_WIDTH-1:0] col_demux_out_data_1;
	wire [DATA_WIDTH-1:0] col_demux_out_data_2;
	wire [DATA_WIDTH-1:0] col_demux_out_data_3;
	wire [DATA_WIDTH-1:0] col_demux_out_data_4;
	wire [DATA_WIDTH-1:0] col_demux_out_data_5;
	wire [DATA_WIDTH-1:0] col_demux_out_data_6;
	wire [DATA_WIDTH-1:0] col_demux_out_data_7;
	wire [DATA_WIDTH-1:0] col_demux_out_data_8;
	wire [DATA_WIDTH-1:0] col_demux_out_data_9;
	wire [DATA_WIDTH-1:0] col_demux_out_data_10;
	wire [DATA_WIDTH-1:0] col_demux_out_data_11;
	wire [DATA_WIDTH-1:0] col_demux_out_data_12;
	wire [DATA_WIDTH-1:0] col_demux_out_data_13;
	wire [DATA_WIDTH-1:0] col_demux_out_data_14;
	wire [DATA_WIDTH-1:0] col_demux_out_data_15;
	wire [DATA_WIDTH-1:0] col_demux_out_data_16;
	wire [DATA_WIDTH-1:0] col_demux_out_data_17;
	wire [DATA_WIDTH-1:0] col_demux_out_data_18;
	wire [DATA_WIDTH-1:0] col_demux_out_data_19;
	wire [DATA_WIDTH-1:0] col_demux_out_data_20;
	wire [DATA_WIDTH-1:0] col_demux_out_data_21;
	wire [DATA_WIDTH-1:0] col_demux_out_data_22;
	wire [DATA_WIDTH-1:0] col_demux_out_data_23;
	wire [DATA_WIDTH-1:0] col_demux_out_data_24;
	wire [DATA_WIDTH-1:0] col_demux_out_data_25;
	wire [DATA_WIDTH-1:0] col_demux_out_data_26;
	wire [DATA_WIDTH-1:0] col_demux_out_data_27;
	wire [DATA_WIDTH-1:0] col_demux_out_data_28;
	wire [DATA_WIDTH-1:0] col_demux_out_data_29;
	wire [DATA_WIDTH-1:0] col_demux_out_data_30;
	wire [DATA_WIDTH-1:0] col_demux_out_data_31;
	demux_1_to_32  col_demux (
		.select (col_select),
		.in_data (in_row),
		.out_data_0 (col_demux_out_data_0),
		.out_data_1 (col_demux_out_data_1),
		.out_data_2 (col_demux_out_data_2),
		.out_data_3 (col_demux_out_data_3),
		.out_data_4 (col_demux_out_data_4),
		.out_data_5 (col_demux_out_data_5),
		.out_data_6 (col_demux_out_data_6),
		.out_data_7 (col_demux_out_data_7),
		.out_data_8 (col_demux_out_data_8),
		.out_data_9 (col_demux_out_data_9),
		.out_data_10 (col_demux_out_data_10),
		.out_data_11 (col_demux_out_data_11),
		.out_data_12 (col_demux_out_data_12),
		.out_data_13 (col_demux_out_data_13),
		.out_data_14 (col_demux_out_data_14),
		.out_data_15 (col_demux_out_data_15),
		.out_data_16 (col_demux_out_data_16),
		.out_data_17 (col_demux_out_data_17),
		.out_data_18 (col_demux_out_data_18),
		.out_data_19 (col_demux_out_data_19),
		.out_data_20 (col_demux_out_data_20),
		.out_data_21 (col_demux_out_data_21),
		.out_data_22 (col_demux_out_data_22),
		.out_data_23 (col_demux_out_data_23),
		.out_data_24 (col_demux_out_data_24),
		.out_data_25 (col_demux_out_data_25),
		.out_data_26 (col_demux_out_data_26),
		.out_data_27 (col_demux_out_data_27),
		.out_data_28 (col_demux_out_data_28),
		.out_data_29 (col_demux_out_data_29),
		.out_data_30 (col_demux_out_data_30),
		.out_data_31 (col_demux_out_data_31)
	);
	////////////////////////////////////////////////////
	// FIFO Instantiations
	////////////////////////////////////////////////////
	wire signed [DATA_WIDTH-1:0] row_fifo_0_out;
	fifo  row_fifo_0 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_0),
		.out_data (row_fifo_0_out),
		.full (row_fifo_0_full),
		.empty(row_fifo_0_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_1_out;
	fifo  row_fifo_1 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_1),
		.out_data (row_fifo_1_out),
		.full (row_fifo_1_full),
		.empty(row_fifo_1_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_2_out;
	fifo  row_fifo_2 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_2),
		.out_data (row_fifo_2_out),
		.full (row_fifo_2_full),
		.empty(row_fifo_2_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_3_out;
	fifo  row_fifo_3 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_3),
		.out_data (row_fifo_3_out),
		.full (row_fifo_3_full),
		.empty(row_fifo_3_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_4_out;
	fifo  row_fifo_4 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_4),
		.out_data (row_fifo_4_out),
		.full (row_fifo_4_full),
		.empty(row_fifo_4_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_5_out;
	fifo  row_fifo_5 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_5),
		.out_data (row_fifo_5_out),
		.full (row_fifo_5_full),
		.empty(row_fifo_5_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_6_out;
	fifo  row_fifo_6 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_6),
		.out_data (row_fifo_6_out),
		.full (row_fifo_6_full),
		.empty(row_fifo_6_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_7_out;
	fifo  row_fifo_7 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_7),
		.out_data (row_fifo_7_out),
		.full (row_fifo_7_full),
		.empty(row_fifo_7_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_8_out;
	fifo  row_fifo_8 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_8),
		.out_data (row_fifo_8_out),
		.full (row_fifo_8_full),
		.empty(row_fifo_8_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_9_out;
	fifo  row_fifo_9 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_9),
		.out_data (row_fifo_9_out),
		.full (row_fifo_9_full),
		.empty(row_fifo_9_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_10_out;
	fifo  row_fifo_10 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_10),
		.out_data (row_fifo_10_out),
		.full (row_fifo_10_full),
		.empty(row_fifo_10_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_11_out;
	fifo  row_fifo_11 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_11),
		.out_data (row_fifo_11_out),
		.full (row_fifo_11_full),
		.empty(row_fifo_11_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_12_out;
	fifo  row_fifo_12 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_12),
		.out_data (row_fifo_12_out),
		.full (row_fifo_12_full),
		.empty(row_fifo_12_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_13_out;
	fifo  row_fifo_13 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_13),
		.out_data (row_fifo_13_out),
		.full (row_fifo_13_full),
		.empty(row_fifo_13_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_14_out;
	fifo  row_fifo_14 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_14),
		.out_data (row_fifo_14_out),
		.full (row_fifo_14_full),
		.empty(row_fifo_14_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_15_out;
	fifo  row_fifo_15 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_15),
		.out_data (row_fifo_15_out),
		.full (row_fifo_15_full),
		.empty(row_fifo_15_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_16_out;
	fifo  row_fifo_16 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_16),
		.out_data (row_fifo_16_out),
		.full (row_fifo_16_full),
		.empty(row_fifo_16_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_17_out;
	fifo  row_fifo_17 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_17),
		.out_data (row_fifo_17_out),
		.full (row_fifo_17_full),
		.empty(row_fifo_17_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_18_out;
	fifo  row_fifo_18 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_18),
		.out_data (row_fifo_18_out),
		.full (row_fifo_18_full),
		.empty(row_fifo_18_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_19_out;
	fifo  row_fifo_19 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_19),
		.out_data (row_fifo_19_out),
		.full (row_fifo_19_full),
		.empty(row_fifo_19_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_20_out;
	fifo  row_fifo_20 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_20),
		.out_data (row_fifo_20_out),
		.full (row_fifo_20_full),
		.empty(row_fifo_20_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_21_out;
	fifo  row_fifo_21 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_21),
		.out_data (row_fifo_21_out),
		.full (row_fifo_21_full),
		.empty(row_fifo_21_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_22_out;
	fifo  row_fifo_22 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_22),
		.out_data (row_fifo_22_out),
		.full (row_fifo_22_full),
		.empty(row_fifo_22_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_23_out;
	fifo  row_fifo_23 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_23),
		.out_data (row_fifo_23_out),
		.full (row_fifo_23_full),
		.empty(row_fifo_23_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_24_out;
	fifo  row_fifo_24 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_24),
		.out_data (row_fifo_24_out),
		.full (row_fifo_24_full),
		.empty(row_fifo_24_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_25_out;
	fifo  row_fifo_25 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_25),
		.out_data (row_fifo_25_out),
		.full (row_fifo_25_full),
		.empty(row_fifo_25_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_26_out;
	fifo  row_fifo_26 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_26),
		.out_data (row_fifo_26_out),
		.full (row_fifo_26_full),
		.empty(row_fifo_26_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_27_out;
	fifo  row_fifo_27 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_27),
		.out_data (row_fifo_27_out),
		.full (row_fifo_27_full),
		.empty(row_fifo_27_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_28_out;
	fifo  row_fifo_28 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_28),
		.out_data (row_fifo_28_out),
		.full (row_fifo_28_full),
		.empty(row_fifo_28_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_29_out;
	fifo  row_fifo_29 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_29),
		.out_data (row_fifo_29_out),
		.full (row_fifo_29_full),
		.empty(row_fifo_29_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_30_out;
	fifo  row_fifo_30 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_30),
		.out_data (row_fifo_30_out),
		.full (row_fifo_30_full),
		.empty(row_fifo_30_empty)
	);
	wire signed [DATA_WIDTH-1:0] row_fifo_31_out;
	fifo  row_fifo_31 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (row_demux_out_data_31),
		.out_data (row_fifo_31_out),
		.full (row_fifo_31_full),
		.empty(row_fifo_31_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_0_out;
	fifo  col_fifo_0 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_0),
		.out_data (col_fifo_0_out),
		.full (col_fifo_0_full),
		.empty(col_fifo_0_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_1_out;
	fifo  col_fifo_1 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_1),
		.out_data (col_fifo_1_out),
		.full (col_fifo_1_full),
		.empty(col_fifo_1_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_2_out;
	fifo  col_fifo_2 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_2),
		.out_data (col_fifo_2_out),
		.full (col_fifo_2_full),
		.empty(col_fifo_2_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_3_out;
	fifo  col_fifo_3 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_3),
		.out_data (col_fifo_3_out),
		.full (col_fifo_3_full),
		.empty(col_fifo_3_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_4_out;
	fifo  col_fifo_4 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_4),
		.out_data (col_fifo_4_out),
		.full (col_fifo_4_full),
		.empty(col_fifo_4_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_5_out;
	fifo  col_fifo_5 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_5),
		.out_data (col_fifo_5_out),
		.full (col_fifo_5_full),
		.empty(col_fifo_5_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_6_out;
	fifo  col_fifo_6 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_6),
		.out_data (col_fifo_6_out),
		.full (col_fifo_6_full),
		.empty(col_fifo_6_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_7_out;
	fifo  col_fifo_7 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_7),
		.out_data (col_fifo_7_out),
		.full (col_fifo_7_full),
		.empty(col_fifo_7_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_8_out;
	fifo  col_fifo_8 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_8),
		.out_data (col_fifo_8_out),
		.full (col_fifo_8_full),
		.empty(col_fifo_8_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_9_out;
	fifo  col_fifo_9 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_9),
		.out_data (col_fifo_9_out),
		.full (col_fifo_9_full),
		.empty(col_fifo_9_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_10_out;
	fifo  col_fifo_10 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_10),
		.out_data (col_fifo_10_out),
		.full (col_fifo_10_full),
		.empty(col_fifo_10_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_11_out;
	fifo  col_fifo_11 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_11),
		.out_data (col_fifo_11_out),
		.full (col_fifo_11_full),
		.empty(col_fifo_11_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_12_out;
	fifo  col_fifo_12 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_12),
		.out_data (col_fifo_12_out),
		.full (col_fifo_12_full),
		.empty(col_fifo_12_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_13_out;
	fifo  col_fifo_13 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_13),
		.out_data (col_fifo_13_out),
		.full (col_fifo_13_full),
		.empty(col_fifo_13_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_14_out;
	fifo  col_fifo_14 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_14),
		.out_data (col_fifo_14_out),
		.full (col_fifo_14_full),
		.empty(col_fifo_14_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_15_out;
	fifo  col_fifo_15 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_15),
		.out_data (col_fifo_15_out),
		.full (col_fifo_15_full),
		.empty(col_fifo_15_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_16_out;
	fifo  col_fifo_16 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_16),
		.out_data (col_fifo_16_out),
		.full (col_fifo_16_full),
		.empty(col_fifo_16_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_17_out;
	fifo  col_fifo_17 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_17),
		.out_data (col_fifo_17_out),
		.full (col_fifo_17_full),
		.empty(col_fifo_17_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_18_out;
	fifo  col_fifo_18 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_18),
		.out_data (col_fifo_18_out),
		.full (col_fifo_18_full),
		.empty(col_fifo_18_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_19_out;
	fifo  col_fifo_19 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_19),
		.out_data (col_fifo_19_out),
		.full (col_fifo_19_full),
		.empty(col_fifo_19_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_20_out;
	fifo  col_fifo_20 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_20),
		.out_data (col_fifo_20_out),
		.full (col_fifo_20_full),
		.empty(col_fifo_20_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_21_out;
	fifo  col_fifo_21 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_21),
		.out_data (col_fifo_21_out),
		.full (col_fifo_21_full),
		.empty(col_fifo_21_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_22_out;
	fifo  col_fifo_22 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_22),
		.out_data (col_fifo_22_out),
		.full (col_fifo_22_full),
		.empty(col_fifo_22_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_23_out;
	fifo  col_fifo_23 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_23),
		.out_data (col_fifo_23_out),
		.full (col_fifo_23_full),
		.empty(col_fifo_23_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_24_out;
	fifo  col_fifo_24 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_24),
		.out_data (col_fifo_24_out),
		.full (col_fifo_24_full),
		.empty(col_fifo_24_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_25_out;
	fifo  col_fifo_25 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_25),
		.out_data (col_fifo_25_out),
		.full (col_fifo_25_full),
		.empty(col_fifo_25_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_26_out;
	fifo  col_fifo_26 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_26),
		.out_data (col_fifo_26_out),
		.full (col_fifo_26_full),
		.empty(col_fifo_26_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_27_out;
	fifo  col_fifo_27 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_27),
		.out_data (col_fifo_27_out),
		.full (col_fifo_27_full),
		.empty(col_fifo_27_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_28_out;
	fifo  col_fifo_28 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_28),
		.out_data (col_fifo_28_out),
		.full (col_fifo_28_full),
		.empty(col_fifo_28_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_29_out;
	fifo  col_fifo_29 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_29),
		.out_data (col_fifo_29_out),
		.full (col_fifo_29_full),
		.empty(col_fifo_29_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_30_out;
	fifo  col_fifo_30 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_30),
		.out_data (col_fifo_30_out),
		.full (col_fifo_30_full),
		.empty(col_fifo_30_empty)
	);
	wire signed [DATA_WIDTH-1:0] col_fifo_31_out;
	fifo  col_fifo_31 (
		.clk (clk),
		.rstn (rstn),
		.w_en (w_en),
		.r_en (r_en),
		.in_data (col_demux_out_data_31),
		.out_data (col_fifo_31_out),
		.full (col_fifo_31_full),
		.empty(col_fifo_31_empty)
	);
	////////////////////////////////////////////////////
	// MAC PE Instantiations
	////////////////////////////////////////////////////
	wire signed [DATA_WIDTH-1:0] out_row_0_0;
	wire signed [DATA_WIDTH-1:0] out_col_0_0;
	wire signed [DATA_WIDTH-1:0] out_data_0_0;
	integer_mac_pe mac_pe_0_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_0_out),
		.in_col (col_fifo_0_out),
		.out_row (out_row_0_0),
		.out_col (out_col_0_0),
		.out_data (out_data_0_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_1;
	wire signed [DATA_WIDTH-1:0] out_col_0_1;
	wire signed [DATA_WIDTH-1:0] out_data_0_1;
	integer_mac_pe mac_pe_0_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_0),
		.in_col (col_fifo_1_out),
		.out_row (out_row_0_1),
		.out_col (out_col_0_1),
		.out_data (out_data_0_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_2;
	wire signed [DATA_WIDTH-1:0] out_col_0_2;
	wire signed [DATA_WIDTH-1:0] out_data_0_2;
	integer_mac_pe mac_pe_0_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_1),
		.in_col (col_fifo_2_out),
		.out_row (out_row_0_2),
		.out_col (out_col_0_2),
		.out_data (out_data_0_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_3;
	wire signed [DATA_WIDTH-1:0] out_col_0_3;
	wire signed [DATA_WIDTH-1:0] out_data_0_3;
	integer_mac_pe mac_pe_0_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_2),
		.in_col (col_fifo_3_out),
		.out_row (out_row_0_3),
		.out_col (out_col_0_3),
		.out_data (out_data_0_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_4;
	wire signed [DATA_WIDTH-1:0] out_col_0_4;
	wire signed [DATA_WIDTH-1:0] out_data_0_4;
	integer_mac_pe mac_pe_0_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_3),
		.in_col (col_fifo_4_out),
		.out_row (out_row_0_4),
		.out_col (out_col_0_4),
		.out_data (out_data_0_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_5;
	wire signed [DATA_WIDTH-1:0] out_col_0_5;
	wire signed [DATA_WIDTH-1:0] out_data_0_5;
	integer_mac_pe mac_pe_0_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_4),
		.in_col (col_fifo_5_out),
		.out_row (out_row_0_5),
		.out_col (out_col_0_5),
		.out_data (out_data_0_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_6;
	wire signed [DATA_WIDTH-1:0] out_col_0_6;
	wire signed [DATA_WIDTH-1:0] out_data_0_6;
	integer_mac_pe mac_pe_0_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_5),
		.in_col (col_fifo_6_out),
		.out_row (out_row_0_6),
		.out_col (out_col_0_6),
		.out_data (out_data_0_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_7;
	wire signed [DATA_WIDTH-1:0] out_col_0_7;
	wire signed [DATA_WIDTH-1:0] out_data_0_7;
	integer_mac_pe mac_pe_0_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_6),
		.in_col (col_fifo_7_out),
		.out_row (out_row_0_7),
		.out_col (out_col_0_7),
		.out_data (out_data_0_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_8;
	wire signed [DATA_WIDTH-1:0] out_col_0_8;
	wire signed [DATA_WIDTH-1:0] out_data_0_8;
	integer_mac_pe mac_pe_0_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_7),
		.in_col (col_fifo_8_out),
		.out_row (out_row_0_8),
		.out_col (out_col_0_8),
		.out_data (out_data_0_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_9;
	wire signed [DATA_WIDTH-1:0] out_col_0_9;
	wire signed [DATA_WIDTH-1:0] out_data_0_9;
	integer_mac_pe mac_pe_0_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_8),
		.in_col (col_fifo_9_out),
		.out_row (out_row_0_9),
		.out_col (out_col_0_9),
		.out_data (out_data_0_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_10;
	wire signed [DATA_WIDTH-1:0] out_col_0_10;
	wire signed [DATA_WIDTH-1:0] out_data_0_10;
	integer_mac_pe mac_pe_0_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_9),
		.in_col (col_fifo_10_out),
		.out_row (out_row_0_10),
		.out_col (out_col_0_10),
		.out_data (out_data_0_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_11;
	wire signed [DATA_WIDTH-1:0] out_col_0_11;
	wire signed [DATA_WIDTH-1:0] out_data_0_11;
	integer_mac_pe mac_pe_0_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_10),
		.in_col (col_fifo_11_out),
		.out_row (out_row_0_11),
		.out_col (out_col_0_11),
		.out_data (out_data_0_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_12;
	wire signed [DATA_WIDTH-1:0] out_col_0_12;
	wire signed [DATA_WIDTH-1:0] out_data_0_12;
	integer_mac_pe mac_pe_0_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_11),
		.in_col (col_fifo_12_out),
		.out_row (out_row_0_12),
		.out_col (out_col_0_12),
		.out_data (out_data_0_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_13;
	wire signed [DATA_WIDTH-1:0] out_col_0_13;
	wire signed [DATA_WIDTH-1:0] out_data_0_13;
	integer_mac_pe mac_pe_0_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_12),
		.in_col (col_fifo_13_out),
		.out_row (out_row_0_13),
		.out_col (out_col_0_13),
		.out_data (out_data_0_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_14;
	wire signed [DATA_WIDTH-1:0] out_col_0_14;
	wire signed [DATA_WIDTH-1:0] out_data_0_14;
	integer_mac_pe mac_pe_0_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_13),
		.in_col (col_fifo_14_out),
		.out_row (out_row_0_14),
		.out_col (out_col_0_14),
		.out_data (out_data_0_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_15;
	wire signed [DATA_WIDTH-1:0] out_col_0_15;
	wire signed [DATA_WIDTH-1:0] out_data_0_15;
	integer_mac_pe mac_pe_0_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_14),
		.in_col (col_fifo_15_out),
		.out_row (out_row_0_15),
		.out_col (out_col_0_15),
		.out_data (out_data_0_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_16;
	wire signed [DATA_WIDTH-1:0] out_col_0_16;
	wire signed [DATA_WIDTH-1:0] out_data_0_16;
	integer_mac_pe mac_pe_0_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_15),
		.in_col (col_fifo_16_out),
		.out_row (out_row_0_16),
		.out_col (out_col_0_16),
		.out_data (out_data_0_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_17;
	wire signed [DATA_WIDTH-1:0] out_col_0_17;
	wire signed [DATA_WIDTH-1:0] out_data_0_17;
	integer_mac_pe mac_pe_0_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_16),
		.in_col (col_fifo_17_out),
		.out_row (out_row_0_17),
		.out_col (out_col_0_17),
		.out_data (out_data_0_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_18;
	wire signed [DATA_WIDTH-1:0] out_col_0_18;
	wire signed [DATA_WIDTH-1:0] out_data_0_18;
	integer_mac_pe mac_pe_0_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_17),
		.in_col (col_fifo_18_out),
		.out_row (out_row_0_18),
		.out_col (out_col_0_18),
		.out_data (out_data_0_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_19;
	wire signed [DATA_WIDTH-1:0] out_col_0_19;
	wire signed [DATA_WIDTH-1:0] out_data_0_19;
	integer_mac_pe mac_pe_0_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_18),
		.in_col (col_fifo_19_out),
		.out_row (out_row_0_19),
		.out_col (out_col_0_19),
		.out_data (out_data_0_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_20;
	wire signed [DATA_WIDTH-1:0] out_col_0_20;
	wire signed [DATA_WIDTH-1:0] out_data_0_20;
	integer_mac_pe mac_pe_0_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_19),
		.in_col (col_fifo_20_out),
		.out_row (out_row_0_20),
		.out_col (out_col_0_20),
		.out_data (out_data_0_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_21;
	wire signed [DATA_WIDTH-1:0] out_col_0_21;
	wire signed [DATA_WIDTH-1:0] out_data_0_21;
	integer_mac_pe mac_pe_0_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_20),
		.in_col (col_fifo_21_out),
		.out_row (out_row_0_21),
		.out_col (out_col_0_21),
		.out_data (out_data_0_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_22;
	wire signed [DATA_WIDTH-1:0] out_col_0_22;
	wire signed [DATA_WIDTH-1:0] out_data_0_22;
	integer_mac_pe mac_pe_0_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_21),
		.in_col (col_fifo_22_out),
		.out_row (out_row_0_22),
		.out_col (out_col_0_22),
		.out_data (out_data_0_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_23;
	wire signed [DATA_WIDTH-1:0] out_col_0_23;
	wire signed [DATA_WIDTH-1:0] out_data_0_23;
	integer_mac_pe mac_pe_0_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_22),
		.in_col (col_fifo_23_out),
		.out_row (out_row_0_23),
		.out_col (out_col_0_23),
		.out_data (out_data_0_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_24;
	wire signed [DATA_WIDTH-1:0] out_col_0_24;
	wire signed [DATA_WIDTH-1:0] out_data_0_24;
	integer_mac_pe mac_pe_0_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_23),
		.in_col (col_fifo_24_out),
		.out_row (out_row_0_24),
		.out_col (out_col_0_24),
		.out_data (out_data_0_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_25;
	wire signed [DATA_WIDTH-1:0] out_col_0_25;
	wire signed [DATA_WIDTH-1:0] out_data_0_25;
	integer_mac_pe mac_pe_0_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_24),
		.in_col (col_fifo_25_out),
		.out_row (out_row_0_25),
		.out_col (out_col_0_25),
		.out_data (out_data_0_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_26;
	wire signed [DATA_WIDTH-1:0] out_col_0_26;
	wire signed [DATA_WIDTH-1:0] out_data_0_26;
	integer_mac_pe mac_pe_0_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_25),
		.in_col (col_fifo_26_out),
		.out_row (out_row_0_26),
		.out_col (out_col_0_26),
		.out_data (out_data_0_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_27;
	wire signed [DATA_WIDTH-1:0] out_col_0_27;
	wire signed [DATA_WIDTH-1:0] out_data_0_27;
	integer_mac_pe mac_pe_0_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_26),
		.in_col (col_fifo_27_out),
		.out_row (out_row_0_27),
		.out_col (out_col_0_27),
		.out_data (out_data_0_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_28;
	wire signed [DATA_WIDTH-1:0] out_col_0_28;
	wire signed [DATA_WIDTH-1:0] out_data_0_28;
	integer_mac_pe mac_pe_0_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_27),
		.in_col (col_fifo_28_out),
		.out_row (out_row_0_28),
		.out_col (out_col_0_28),
		.out_data (out_data_0_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_29;
	wire signed [DATA_WIDTH-1:0] out_col_0_29;
	wire signed [DATA_WIDTH-1:0] out_data_0_29;
	integer_mac_pe mac_pe_0_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_28),
		.in_col (col_fifo_29_out),
		.out_row (out_row_0_29),
		.out_col (out_col_0_29),
		.out_data (out_data_0_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_30;
	wire signed [DATA_WIDTH-1:0] out_col_0_30;
	wire signed [DATA_WIDTH-1:0] out_data_0_30;
	integer_mac_pe mac_pe_0_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_29),
		.in_col (col_fifo_30_out),
		.out_row (out_row_0_30),
		.out_col (out_col_0_30),
		.out_data (out_data_0_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_0_31;
	wire signed [DATA_WIDTH-1:0] out_col_0_31;
	wire signed [DATA_WIDTH-1:0] out_data_0_31;
	integer_mac_pe mac_pe_0_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_0_30),
		.in_col (col_fifo_31_out),
		.out_row (out_row_0_31),
		.out_col (out_col_0_31),
		.out_data (out_data_0_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_0;
	wire signed [DATA_WIDTH-1:0] out_col_1_0;
	wire signed [DATA_WIDTH-1:0] out_data_1_0;
	integer_mac_pe mac_pe_1_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_1_out),
		.in_col (out_col_0_0),
		.out_row (out_row_1_0),
		.out_col (out_col_1_0),
		.out_data (out_data_1_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_1;
	wire signed [DATA_WIDTH-1:0] out_col_1_1;
	wire signed [DATA_WIDTH-1:0] out_data_1_1;
	integer_mac_pe mac_pe_1_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_0),
		.in_col (out_col_0_1),
		.out_row (out_row_1_1),
		.out_col (out_col_1_1),
		.out_data (out_data_1_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_2;
	wire signed [DATA_WIDTH-1:0] out_col_1_2;
	wire signed [DATA_WIDTH-1:0] out_data_1_2;
	integer_mac_pe mac_pe_1_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_1),
		.in_col (out_col_0_2),
		.out_row (out_row_1_2),
		.out_col (out_col_1_2),
		.out_data (out_data_1_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_3;
	wire signed [DATA_WIDTH-1:0] out_col_1_3;
	wire signed [DATA_WIDTH-1:0] out_data_1_3;
	integer_mac_pe mac_pe_1_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_2),
		.in_col (out_col_0_3),
		.out_row (out_row_1_3),
		.out_col (out_col_1_3),
		.out_data (out_data_1_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_4;
	wire signed [DATA_WIDTH-1:0] out_col_1_4;
	wire signed [DATA_WIDTH-1:0] out_data_1_4;
	integer_mac_pe mac_pe_1_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_3),
		.in_col (out_col_0_4),
		.out_row (out_row_1_4),
		.out_col (out_col_1_4),
		.out_data (out_data_1_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_5;
	wire signed [DATA_WIDTH-1:0] out_col_1_5;
	wire signed [DATA_WIDTH-1:0] out_data_1_5;
	integer_mac_pe mac_pe_1_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_4),
		.in_col (out_col_0_5),
		.out_row (out_row_1_5),
		.out_col (out_col_1_5),
		.out_data (out_data_1_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_6;
	wire signed [DATA_WIDTH-1:0] out_col_1_6;
	wire signed [DATA_WIDTH-1:0] out_data_1_6;
	integer_mac_pe mac_pe_1_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_5),
		.in_col (out_col_0_6),
		.out_row (out_row_1_6),
		.out_col (out_col_1_6),
		.out_data (out_data_1_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_7;
	wire signed [DATA_WIDTH-1:0] out_col_1_7;
	wire signed [DATA_WIDTH-1:0] out_data_1_7;
	integer_mac_pe mac_pe_1_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_6),
		.in_col (out_col_0_7),
		.out_row (out_row_1_7),
		.out_col (out_col_1_7),
		.out_data (out_data_1_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_8;
	wire signed [DATA_WIDTH-1:0] out_col_1_8;
	wire signed [DATA_WIDTH-1:0] out_data_1_8;
	integer_mac_pe mac_pe_1_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_7),
		.in_col (out_col_0_8),
		.out_row (out_row_1_8),
		.out_col (out_col_1_8),
		.out_data (out_data_1_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_9;
	wire signed [DATA_WIDTH-1:0] out_col_1_9;
	wire signed [DATA_WIDTH-1:0] out_data_1_9;
	integer_mac_pe mac_pe_1_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_8),
		.in_col (out_col_0_9),
		.out_row (out_row_1_9),
		.out_col (out_col_1_9),
		.out_data (out_data_1_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_10;
	wire signed [DATA_WIDTH-1:0] out_col_1_10;
	wire signed [DATA_WIDTH-1:0] out_data_1_10;
	integer_mac_pe mac_pe_1_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_9),
		.in_col (out_col_0_10),
		.out_row (out_row_1_10),
		.out_col (out_col_1_10),
		.out_data (out_data_1_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_11;
	wire signed [DATA_WIDTH-1:0] out_col_1_11;
	wire signed [DATA_WIDTH-1:0] out_data_1_11;
	integer_mac_pe mac_pe_1_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_10),
		.in_col (out_col_0_11),
		.out_row (out_row_1_11),
		.out_col (out_col_1_11),
		.out_data (out_data_1_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_12;
	wire signed [DATA_WIDTH-1:0] out_col_1_12;
	wire signed [DATA_WIDTH-1:0] out_data_1_12;
	integer_mac_pe mac_pe_1_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_11),
		.in_col (out_col_0_12),
		.out_row (out_row_1_12),
		.out_col (out_col_1_12),
		.out_data (out_data_1_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_13;
	wire signed [DATA_WIDTH-1:0] out_col_1_13;
	wire signed [DATA_WIDTH-1:0] out_data_1_13;
	integer_mac_pe mac_pe_1_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_12),
		.in_col (out_col_0_13),
		.out_row (out_row_1_13),
		.out_col (out_col_1_13),
		.out_data (out_data_1_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_14;
	wire signed [DATA_WIDTH-1:0] out_col_1_14;
	wire signed [DATA_WIDTH-1:0] out_data_1_14;
	integer_mac_pe mac_pe_1_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_13),
		.in_col (out_col_0_14),
		.out_row (out_row_1_14),
		.out_col (out_col_1_14),
		.out_data (out_data_1_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_15;
	wire signed [DATA_WIDTH-1:0] out_col_1_15;
	wire signed [DATA_WIDTH-1:0] out_data_1_15;
	integer_mac_pe mac_pe_1_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_14),
		.in_col (out_col_0_15),
		.out_row (out_row_1_15),
		.out_col (out_col_1_15),
		.out_data (out_data_1_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_16;
	wire signed [DATA_WIDTH-1:0] out_col_1_16;
	wire signed [DATA_WIDTH-1:0] out_data_1_16;
	integer_mac_pe mac_pe_1_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_15),
		.in_col (out_col_0_16),
		.out_row (out_row_1_16),
		.out_col (out_col_1_16),
		.out_data (out_data_1_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_17;
	wire signed [DATA_WIDTH-1:0] out_col_1_17;
	wire signed [DATA_WIDTH-1:0] out_data_1_17;
	integer_mac_pe mac_pe_1_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_16),
		.in_col (out_col_0_17),
		.out_row (out_row_1_17),
		.out_col (out_col_1_17),
		.out_data (out_data_1_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_18;
	wire signed [DATA_WIDTH-1:0] out_col_1_18;
	wire signed [DATA_WIDTH-1:0] out_data_1_18;
	integer_mac_pe mac_pe_1_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_17),
		.in_col (out_col_0_18),
		.out_row (out_row_1_18),
		.out_col (out_col_1_18),
		.out_data (out_data_1_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_19;
	wire signed [DATA_WIDTH-1:0] out_col_1_19;
	wire signed [DATA_WIDTH-1:0] out_data_1_19;
	integer_mac_pe mac_pe_1_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_18),
		.in_col (out_col_0_19),
		.out_row (out_row_1_19),
		.out_col (out_col_1_19),
		.out_data (out_data_1_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_20;
	wire signed [DATA_WIDTH-1:0] out_col_1_20;
	wire signed [DATA_WIDTH-1:0] out_data_1_20;
	integer_mac_pe mac_pe_1_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_19),
		.in_col (out_col_0_20),
		.out_row (out_row_1_20),
		.out_col (out_col_1_20),
		.out_data (out_data_1_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_21;
	wire signed [DATA_WIDTH-1:0] out_col_1_21;
	wire signed [DATA_WIDTH-1:0] out_data_1_21;
	integer_mac_pe mac_pe_1_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_20),
		.in_col (out_col_0_21),
		.out_row (out_row_1_21),
		.out_col (out_col_1_21),
		.out_data (out_data_1_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_22;
	wire signed [DATA_WIDTH-1:0] out_col_1_22;
	wire signed [DATA_WIDTH-1:0] out_data_1_22;
	integer_mac_pe mac_pe_1_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_21),
		.in_col (out_col_0_22),
		.out_row (out_row_1_22),
		.out_col (out_col_1_22),
		.out_data (out_data_1_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_23;
	wire signed [DATA_WIDTH-1:0] out_col_1_23;
	wire signed [DATA_WIDTH-1:0] out_data_1_23;
	integer_mac_pe mac_pe_1_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_22),
		.in_col (out_col_0_23),
		.out_row (out_row_1_23),
		.out_col (out_col_1_23),
		.out_data (out_data_1_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_24;
	wire signed [DATA_WIDTH-1:0] out_col_1_24;
	wire signed [DATA_WIDTH-1:0] out_data_1_24;
	integer_mac_pe mac_pe_1_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_23),
		.in_col (out_col_0_24),
		.out_row (out_row_1_24),
		.out_col (out_col_1_24),
		.out_data (out_data_1_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_25;
	wire signed [DATA_WIDTH-1:0] out_col_1_25;
	wire signed [DATA_WIDTH-1:0] out_data_1_25;
	integer_mac_pe mac_pe_1_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_24),
		.in_col (out_col_0_25),
		.out_row (out_row_1_25),
		.out_col (out_col_1_25),
		.out_data (out_data_1_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_26;
	wire signed [DATA_WIDTH-1:0] out_col_1_26;
	wire signed [DATA_WIDTH-1:0] out_data_1_26;
	integer_mac_pe mac_pe_1_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_25),
		.in_col (out_col_0_26),
		.out_row (out_row_1_26),
		.out_col (out_col_1_26),
		.out_data (out_data_1_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_27;
	wire signed [DATA_WIDTH-1:0] out_col_1_27;
	wire signed [DATA_WIDTH-1:0] out_data_1_27;
	integer_mac_pe mac_pe_1_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_26),
		.in_col (out_col_0_27),
		.out_row (out_row_1_27),
		.out_col (out_col_1_27),
		.out_data (out_data_1_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_28;
	wire signed [DATA_WIDTH-1:0] out_col_1_28;
	wire signed [DATA_WIDTH-1:0] out_data_1_28;
	integer_mac_pe mac_pe_1_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_27),
		.in_col (out_col_0_28),
		.out_row (out_row_1_28),
		.out_col (out_col_1_28),
		.out_data (out_data_1_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_29;
	wire signed [DATA_WIDTH-1:0] out_col_1_29;
	wire signed [DATA_WIDTH-1:0] out_data_1_29;
	integer_mac_pe mac_pe_1_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_28),
		.in_col (out_col_0_29),
		.out_row (out_row_1_29),
		.out_col (out_col_1_29),
		.out_data (out_data_1_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_30;
	wire signed [DATA_WIDTH-1:0] out_col_1_30;
	wire signed [DATA_WIDTH-1:0] out_data_1_30;
	integer_mac_pe mac_pe_1_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_29),
		.in_col (out_col_0_30),
		.out_row (out_row_1_30),
		.out_col (out_col_1_30),
		.out_data (out_data_1_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_1_31;
	wire signed [DATA_WIDTH-1:0] out_col_1_31;
	wire signed [DATA_WIDTH-1:0] out_data_1_31;
	integer_mac_pe mac_pe_1_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_1_30),
		.in_col (out_col_0_31),
		.out_row (out_row_1_31),
		.out_col (out_col_1_31),
		.out_data (out_data_1_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_0;
	wire signed [DATA_WIDTH-1:0] out_col_2_0;
	wire signed [DATA_WIDTH-1:0] out_data_2_0;
	integer_mac_pe mac_pe_2_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_2_out),
		.in_col (out_col_1_0),
		.out_row (out_row_2_0),
		.out_col (out_col_2_0),
		.out_data (out_data_2_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_1;
	wire signed [DATA_WIDTH-1:0] out_col_2_1;
	wire signed [DATA_WIDTH-1:0] out_data_2_1;
	integer_mac_pe mac_pe_2_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_0),
		.in_col (out_col_1_1),
		.out_row (out_row_2_1),
		.out_col (out_col_2_1),
		.out_data (out_data_2_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_2;
	wire signed [DATA_WIDTH-1:0] out_col_2_2;
	wire signed [DATA_WIDTH-1:0] out_data_2_2;
	integer_mac_pe mac_pe_2_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_1),
		.in_col (out_col_1_2),
		.out_row (out_row_2_2),
		.out_col (out_col_2_2),
		.out_data (out_data_2_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_3;
	wire signed [DATA_WIDTH-1:0] out_col_2_3;
	wire signed [DATA_WIDTH-1:0] out_data_2_3;
	integer_mac_pe mac_pe_2_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_2),
		.in_col (out_col_1_3),
		.out_row (out_row_2_3),
		.out_col (out_col_2_3),
		.out_data (out_data_2_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_4;
	wire signed [DATA_WIDTH-1:0] out_col_2_4;
	wire signed [DATA_WIDTH-1:0] out_data_2_4;
	integer_mac_pe mac_pe_2_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_3),
		.in_col (out_col_1_4),
		.out_row (out_row_2_4),
		.out_col (out_col_2_4),
		.out_data (out_data_2_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_5;
	wire signed [DATA_WIDTH-1:0] out_col_2_5;
	wire signed [DATA_WIDTH-1:0] out_data_2_5;
	integer_mac_pe mac_pe_2_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_4),
		.in_col (out_col_1_5),
		.out_row (out_row_2_5),
		.out_col (out_col_2_5),
		.out_data (out_data_2_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_6;
	wire signed [DATA_WIDTH-1:0] out_col_2_6;
	wire signed [DATA_WIDTH-1:0] out_data_2_6;
	integer_mac_pe mac_pe_2_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_5),
		.in_col (out_col_1_6),
		.out_row (out_row_2_6),
		.out_col (out_col_2_6),
		.out_data (out_data_2_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_7;
	wire signed [DATA_WIDTH-1:0] out_col_2_7;
	wire signed [DATA_WIDTH-1:0] out_data_2_7;
	integer_mac_pe mac_pe_2_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_6),
		.in_col (out_col_1_7),
		.out_row (out_row_2_7),
		.out_col (out_col_2_7),
		.out_data (out_data_2_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_8;
	wire signed [DATA_WIDTH-1:0] out_col_2_8;
	wire signed [DATA_WIDTH-1:0] out_data_2_8;
	integer_mac_pe mac_pe_2_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_7),
		.in_col (out_col_1_8),
		.out_row (out_row_2_8),
		.out_col (out_col_2_8),
		.out_data (out_data_2_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_9;
	wire signed [DATA_WIDTH-1:0] out_col_2_9;
	wire signed [DATA_WIDTH-1:0] out_data_2_9;
	integer_mac_pe mac_pe_2_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_8),
		.in_col (out_col_1_9),
		.out_row (out_row_2_9),
		.out_col (out_col_2_9),
		.out_data (out_data_2_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_10;
	wire signed [DATA_WIDTH-1:0] out_col_2_10;
	wire signed [DATA_WIDTH-1:0] out_data_2_10;
	integer_mac_pe mac_pe_2_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_9),
		.in_col (out_col_1_10),
		.out_row (out_row_2_10),
		.out_col (out_col_2_10),
		.out_data (out_data_2_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_11;
	wire signed [DATA_WIDTH-1:0] out_col_2_11;
	wire signed [DATA_WIDTH-1:0] out_data_2_11;
	integer_mac_pe mac_pe_2_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_10),
		.in_col (out_col_1_11),
		.out_row (out_row_2_11),
		.out_col (out_col_2_11),
		.out_data (out_data_2_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_12;
	wire signed [DATA_WIDTH-1:0] out_col_2_12;
	wire signed [DATA_WIDTH-1:0] out_data_2_12;
	integer_mac_pe mac_pe_2_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_11),
		.in_col (out_col_1_12),
		.out_row (out_row_2_12),
		.out_col (out_col_2_12),
		.out_data (out_data_2_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_13;
	wire signed [DATA_WIDTH-1:0] out_col_2_13;
	wire signed [DATA_WIDTH-1:0] out_data_2_13;
	integer_mac_pe mac_pe_2_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_12),
		.in_col (out_col_1_13),
		.out_row (out_row_2_13),
		.out_col (out_col_2_13),
		.out_data (out_data_2_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_14;
	wire signed [DATA_WIDTH-1:0] out_col_2_14;
	wire signed [DATA_WIDTH-1:0] out_data_2_14;
	integer_mac_pe mac_pe_2_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_13),
		.in_col (out_col_1_14),
		.out_row (out_row_2_14),
		.out_col (out_col_2_14),
		.out_data (out_data_2_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_15;
	wire signed [DATA_WIDTH-1:0] out_col_2_15;
	wire signed [DATA_WIDTH-1:0] out_data_2_15;
	integer_mac_pe mac_pe_2_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_14),
		.in_col (out_col_1_15),
		.out_row (out_row_2_15),
		.out_col (out_col_2_15),
		.out_data (out_data_2_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_16;
	wire signed [DATA_WIDTH-1:0] out_col_2_16;
	wire signed [DATA_WIDTH-1:0] out_data_2_16;
	integer_mac_pe mac_pe_2_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_15),
		.in_col (out_col_1_16),
		.out_row (out_row_2_16),
		.out_col (out_col_2_16),
		.out_data (out_data_2_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_17;
	wire signed [DATA_WIDTH-1:0] out_col_2_17;
	wire signed [DATA_WIDTH-1:0] out_data_2_17;
	integer_mac_pe mac_pe_2_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_16),
		.in_col (out_col_1_17),
		.out_row (out_row_2_17),
		.out_col (out_col_2_17),
		.out_data (out_data_2_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_18;
	wire signed [DATA_WIDTH-1:0] out_col_2_18;
	wire signed [DATA_WIDTH-1:0] out_data_2_18;
	integer_mac_pe mac_pe_2_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_17),
		.in_col (out_col_1_18),
		.out_row (out_row_2_18),
		.out_col (out_col_2_18),
		.out_data (out_data_2_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_19;
	wire signed [DATA_WIDTH-1:0] out_col_2_19;
	wire signed [DATA_WIDTH-1:0] out_data_2_19;
	integer_mac_pe mac_pe_2_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_18),
		.in_col (out_col_1_19),
		.out_row (out_row_2_19),
		.out_col (out_col_2_19),
		.out_data (out_data_2_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_20;
	wire signed [DATA_WIDTH-1:0] out_col_2_20;
	wire signed [DATA_WIDTH-1:0] out_data_2_20;
	integer_mac_pe mac_pe_2_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_19),
		.in_col (out_col_1_20),
		.out_row (out_row_2_20),
		.out_col (out_col_2_20),
		.out_data (out_data_2_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_21;
	wire signed [DATA_WIDTH-1:0] out_col_2_21;
	wire signed [DATA_WIDTH-1:0] out_data_2_21;
	integer_mac_pe mac_pe_2_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_20),
		.in_col (out_col_1_21),
		.out_row (out_row_2_21),
		.out_col (out_col_2_21),
		.out_data (out_data_2_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_22;
	wire signed [DATA_WIDTH-1:0] out_col_2_22;
	wire signed [DATA_WIDTH-1:0] out_data_2_22;
	integer_mac_pe mac_pe_2_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_21),
		.in_col (out_col_1_22),
		.out_row (out_row_2_22),
		.out_col (out_col_2_22),
		.out_data (out_data_2_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_23;
	wire signed [DATA_WIDTH-1:0] out_col_2_23;
	wire signed [DATA_WIDTH-1:0] out_data_2_23;
	integer_mac_pe mac_pe_2_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_22),
		.in_col (out_col_1_23),
		.out_row (out_row_2_23),
		.out_col (out_col_2_23),
		.out_data (out_data_2_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_24;
	wire signed [DATA_WIDTH-1:0] out_col_2_24;
	wire signed [DATA_WIDTH-1:0] out_data_2_24;
	integer_mac_pe mac_pe_2_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_23),
		.in_col (out_col_1_24),
		.out_row (out_row_2_24),
		.out_col (out_col_2_24),
		.out_data (out_data_2_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_25;
	wire signed [DATA_WIDTH-1:0] out_col_2_25;
	wire signed [DATA_WIDTH-1:0] out_data_2_25;
	integer_mac_pe mac_pe_2_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_24),
		.in_col (out_col_1_25),
		.out_row (out_row_2_25),
		.out_col (out_col_2_25),
		.out_data (out_data_2_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_26;
	wire signed [DATA_WIDTH-1:0] out_col_2_26;
	wire signed [DATA_WIDTH-1:0] out_data_2_26;
	integer_mac_pe mac_pe_2_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_25),
		.in_col (out_col_1_26),
		.out_row (out_row_2_26),
		.out_col (out_col_2_26),
		.out_data (out_data_2_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_27;
	wire signed [DATA_WIDTH-1:0] out_col_2_27;
	wire signed [DATA_WIDTH-1:0] out_data_2_27;
	integer_mac_pe mac_pe_2_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_26),
		.in_col (out_col_1_27),
		.out_row (out_row_2_27),
		.out_col (out_col_2_27),
		.out_data (out_data_2_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_28;
	wire signed [DATA_WIDTH-1:0] out_col_2_28;
	wire signed [DATA_WIDTH-1:0] out_data_2_28;
	integer_mac_pe mac_pe_2_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_27),
		.in_col (out_col_1_28),
		.out_row (out_row_2_28),
		.out_col (out_col_2_28),
		.out_data (out_data_2_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_29;
	wire signed [DATA_WIDTH-1:0] out_col_2_29;
	wire signed [DATA_WIDTH-1:0] out_data_2_29;
	integer_mac_pe mac_pe_2_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_28),
		.in_col (out_col_1_29),
		.out_row (out_row_2_29),
		.out_col (out_col_2_29),
		.out_data (out_data_2_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_30;
	wire signed [DATA_WIDTH-1:0] out_col_2_30;
	wire signed [DATA_WIDTH-1:0] out_data_2_30;
	integer_mac_pe mac_pe_2_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_29),
		.in_col (out_col_1_30),
		.out_row (out_row_2_30),
		.out_col (out_col_2_30),
		.out_data (out_data_2_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_2_31;
	wire signed [DATA_WIDTH-1:0] out_col_2_31;
	wire signed [DATA_WIDTH-1:0] out_data_2_31;
	integer_mac_pe mac_pe_2_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_2_30),
		.in_col (out_col_1_31),
		.out_row (out_row_2_31),
		.out_col (out_col_2_31),
		.out_data (out_data_2_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_0;
	wire signed [DATA_WIDTH-1:0] out_col_3_0;
	wire signed [DATA_WIDTH-1:0] out_data_3_0;
	integer_mac_pe mac_pe_3_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_3_out),
		.in_col (out_col_2_0),
		.out_row (out_row_3_0),
		.out_col (out_col_3_0),
		.out_data (out_data_3_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_1;
	wire signed [DATA_WIDTH-1:0] out_col_3_1;
	wire signed [DATA_WIDTH-1:0] out_data_3_1;
	integer_mac_pe mac_pe_3_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_0),
		.in_col (out_col_2_1),
		.out_row (out_row_3_1),
		.out_col (out_col_3_1),
		.out_data (out_data_3_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_2;
	wire signed [DATA_WIDTH-1:0] out_col_3_2;
	wire signed [DATA_WIDTH-1:0] out_data_3_2;
	integer_mac_pe mac_pe_3_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_1),
		.in_col (out_col_2_2),
		.out_row (out_row_3_2),
		.out_col (out_col_3_2),
		.out_data (out_data_3_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_3;
	wire signed [DATA_WIDTH-1:0] out_col_3_3;
	wire signed [DATA_WIDTH-1:0] out_data_3_3;
	integer_mac_pe mac_pe_3_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_2),
		.in_col (out_col_2_3),
		.out_row (out_row_3_3),
		.out_col (out_col_3_3),
		.out_data (out_data_3_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_4;
	wire signed [DATA_WIDTH-1:0] out_col_3_4;
	wire signed [DATA_WIDTH-1:0] out_data_3_4;
	integer_mac_pe mac_pe_3_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_3),
		.in_col (out_col_2_4),
		.out_row (out_row_3_4),
		.out_col (out_col_3_4),
		.out_data (out_data_3_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_5;
	wire signed [DATA_WIDTH-1:0] out_col_3_5;
	wire signed [DATA_WIDTH-1:0] out_data_3_5;
	integer_mac_pe mac_pe_3_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_4),
		.in_col (out_col_2_5),
		.out_row (out_row_3_5),
		.out_col (out_col_3_5),
		.out_data (out_data_3_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_6;
	wire signed [DATA_WIDTH-1:0] out_col_3_6;
	wire signed [DATA_WIDTH-1:0] out_data_3_6;
	integer_mac_pe mac_pe_3_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_5),
		.in_col (out_col_2_6),
		.out_row (out_row_3_6),
		.out_col (out_col_3_6),
		.out_data (out_data_3_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_7;
	wire signed [DATA_WIDTH-1:0] out_col_3_7;
	wire signed [DATA_WIDTH-1:0] out_data_3_7;
	integer_mac_pe mac_pe_3_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_6),
		.in_col (out_col_2_7),
		.out_row (out_row_3_7),
		.out_col (out_col_3_7),
		.out_data (out_data_3_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_8;
	wire signed [DATA_WIDTH-1:0] out_col_3_8;
	wire signed [DATA_WIDTH-1:0] out_data_3_8;
	integer_mac_pe mac_pe_3_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_7),
		.in_col (out_col_2_8),
		.out_row (out_row_3_8),
		.out_col (out_col_3_8),
		.out_data (out_data_3_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_9;
	wire signed [DATA_WIDTH-1:0] out_col_3_9;
	wire signed [DATA_WIDTH-1:0] out_data_3_9;
	integer_mac_pe mac_pe_3_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_8),
		.in_col (out_col_2_9),
		.out_row (out_row_3_9),
		.out_col (out_col_3_9),
		.out_data (out_data_3_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_10;
	wire signed [DATA_WIDTH-1:0] out_col_3_10;
	wire signed [DATA_WIDTH-1:0] out_data_3_10;
	integer_mac_pe mac_pe_3_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_9),
		.in_col (out_col_2_10),
		.out_row (out_row_3_10),
		.out_col (out_col_3_10),
		.out_data (out_data_3_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_11;
	wire signed [DATA_WIDTH-1:0] out_col_3_11;
	wire signed [DATA_WIDTH-1:0] out_data_3_11;
	integer_mac_pe mac_pe_3_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_10),
		.in_col (out_col_2_11),
		.out_row (out_row_3_11),
		.out_col (out_col_3_11),
		.out_data (out_data_3_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_12;
	wire signed [DATA_WIDTH-1:0] out_col_3_12;
	wire signed [DATA_WIDTH-1:0] out_data_3_12;
	integer_mac_pe mac_pe_3_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_11),
		.in_col (out_col_2_12),
		.out_row (out_row_3_12),
		.out_col (out_col_3_12),
		.out_data (out_data_3_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_13;
	wire signed [DATA_WIDTH-1:0] out_col_3_13;
	wire signed [DATA_WIDTH-1:0] out_data_3_13;
	integer_mac_pe mac_pe_3_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_12),
		.in_col (out_col_2_13),
		.out_row (out_row_3_13),
		.out_col (out_col_3_13),
		.out_data (out_data_3_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_14;
	wire signed [DATA_WIDTH-1:0] out_col_3_14;
	wire signed [DATA_WIDTH-1:0] out_data_3_14;
	integer_mac_pe mac_pe_3_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_13),
		.in_col (out_col_2_14),
		.out_row (out_row_3_14),
		.out_col (out_col_3_14),
		.out_data (out_data_3_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_15;
	wire signed [DATA_WIDTH-1:0] out_col_3_15;
	wire signed [DATA_WIDTH-1:0] out_data_3_15;
	integer_mac_pe mac_pe_3_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_14),
		.in_col (out_col_2_15),
		.out_row (out_row_3_15),
		.out_col (out_col_3_15),
		.out_data (out_data_3_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_16;
	wire signed [DATA_WIDTH-1:0] out_col_3_16;
	wire signed [DATA_WIDTH-1:0] out_data_3_16;
	integer_mac_pe mac_pe_3_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_15),
		.in_col (out_col_2_16),
		.out_row (out_row_3_16),
		.out_col (out_col_3_16),
		.out_data (out_data_3_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_17;
	wire signed [DATA_WIDTH-1:0] out_col_3_17;
	wire signed [DATA_WIDTH-1:0] out_data_3_17;
	integer_mac_pe mac_pe_3_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_16),
		.in_col (out_col_2_17),
		.out_row (out_row_3_17),
		.out_col (out_col_3_17),
		.out_data (out_data_3_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_18;
	wire signed [DATA_WIDTH-1:0] out_col_3_18;
	wire signed [DATA_WIDTH-1:0] out_data_3_18;
	integer_mac_pe mac_pe_3_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_17),
		.in_col (out_col_2_18),
		.out_row (out_row_3_18),
		.out_col (out_col_3_18),
		.out_data (out_data_3_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_19;
	wire signed [DATA_WIDTH-1:0] out_col_3_19;
	wire signed [DATA_WIDTH-1:0] out_data_3_19;
	integer_mac_pe mac_pe_3_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_18),
		.in_col (out_col_2_19),
		.out_row (out_row_3_19),
		.out_col (out_col_3_19),
		.out_data (out_data_3_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_20;
	wire signed [DATA_WIDTH-1:0] out_col_3_20;
	wire signed [DATA_WIDTH-1:0] out_data_3_20;
	integer_mac_pe mac_pe_3_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_19),
		.in_col (out_col_2_20),
		.out_row (out_row_3_20),
		.out_col (out_col_3_20),
		.out_data (out_data_3_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_21;
	wire signed [DATA_WIDTH-1:0] out_col_3_21;
	wire signed [DATA_WIDTH-1:0] out_data_3_21;
	integer_mac_pe mac_pe_3_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_20),
		.in_col (out_col_2_21),
		.out_row (out_row_3_21),
		.out_col (out_col_3_21),
		.out_data (out_data_3_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_22;
	wire signed [DATA_WIDTH-1:0] out_col_3_22;
	wire signed [DATA_WIDTH-1:0] out_data_3_22;
	integer_mac_pe mac_pe_3_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_21),
		.in_col (out_col_2_22),
		.out_row (out_row_3_22),
		.out_col (out_col_3_22),
		.out_data (out_data_3_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_23;
	wire signed [DATA_WIDTH-1:0] out_col_3_23;
	wire signed [DATA_WIDTH-1:0] out_data_3_23;
	integer_mac_pe mac_pe_3_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_22),
		.in_col (out_col_2_23),
		.out_row (out_row_3_23),
		.out_col (out_col_3_23),
		.out_data (out_data_3_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_24;
	wire signed [DATA_WIDTH-1:0] out_col_3_24;
	wire signed [DATA_WIDTH-1:0] out_data_3_24;
	integer_mac_pe mac_pe_3_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_23),
		.in_col (out_col_2_24),
		.out_row (out_row_3_24),
		.out_col (out_col_3_24),
		.out_data (out_data_3_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_25;
	wire signed [DATA_WIDTH-1:0] out_col_3_25;
	wire signed [DATA_WIDTH-1:0] out_data_3_25;
	integer_mac_pe mac_pe_3_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_24),
		.in_col (out_col_2_25),
		.out_row (out_row_3_25),
		.out_col (out_col_3_25),
		.out_data (out_data_3_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_26;
	wire signed [DATA_WIDTH-1:0] out_col_3_26;
	wire signed [DATA_WIDTH-1:0] out_data_3_26;
	integer_mac_pe mac_pe_3_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_25),
		.in_col (out_col_2_26),
		.out_row (out_row_3_26),
		.out_col (out_col_3_26),
		.out_data (out_data_3_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_27;
	wire signed [DATA_WIDTH-1:0] out_col_3_27;
	wire signed [DATA_WIDTH-1:0] out_data_3_27;
	integer_mac_pe mac_pe_3_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_26),
		.in_col (out_col_2_27),
		.out_row (out_row_3_27),
		.out_col (out_col_3_27),
		.out_data (out_data_3_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_28;
	wire signed [DATA_WIDTH-1:0] out_col_3_28;
	wire signed [DATA_WIDTH-1:0] out_data_3_28;
	integer_mac_pe mac_pe_3_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_27),
		.in_col (out_col_2_28),
		.out_row (out_row_3_28),
		.out_col (out_col_3_28),
		.out_data (out_data_3_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_29;
	wire signed [DATA_WIDTH-1:0] out_col_3_29;
	wire signed [DATA_WIDTH-1:0] out_data_3_29;
	integer_mac_pe mac_pe_3_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_28),
		.in_col (out_col_2_29),
		.out_row (out_row_3_29),
		.out_col (out_col_3_29),
		.out_data (out_data_3_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_30;
	wire signed [DATA_WIDTH-1:0] out_col_3_30;
	wire signed [DATA_WIDTH-1:0] out_data_3_30;
	integer_mac_pe mac_pe_3_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_29),
		.in_col (out_col_2_30),
		.out_row (out_row_3_30),
		.out_col (out_col_3_30),
		.out_data (out_data_3_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_3_31;
	wire signed [DATA_WIDTH-1:0] out_col_3_31;
	wire signed [DATA_WIDTH-1:0] out_data_3_31;
	integer_mac_pe mac_pe_3_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_3_30),
		.in_col (out_col_2_31),
		.out_row (out_row_3_31),
		.out_col (out_col_3_31),
		.out_data (out_data_3_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_0;
	wire signed [DATA_WIDTH-1:0] out_col_4_0;
	wire signed [DATA_WIDTH-1:0] out_data_4_0;
	integer_mac_pe mac_pe_4_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_4_out),
		.in_col (out_col_3_0),
		.out_row (out_row_4_0),
		.out_col (out_col_4_0),
		.out_data (out_data_4_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_1;
	wire signed [DATA_WIDTH-1:0] out_col_4_1;
	wire signed [DATA_WIDTH-1:0] out_data_4_1;
	integer_mac_pe mac_pe_4_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_0),
		.in_col (out_col_3_1),
		.out_row (out_row_4_1),
		.out_col (out_col_4_1),
		.out_data (out_data_4_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_2;
	wire signed [DATA_WIDTH-1:0] out_col_4_2;
	wire signed [DATA_WIDTH-1:0] out_data_4_2;
	integer_mac_pe mac_pe_4_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_1),
		.in_col (out_col_3_2),
		.out_row (out_row_4_2),
		.out_col (out_col_4_2),
		.out_data (out_data_4_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_3;
	wire signed [DATA_WIDTH-1:0] out_col_4_3;
	wire signed [DATA_WIDTH-1:0] out_data_4_3;
	integer_mac_pe mac_pe_4_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_2),
		.in_col (out_col_3_3),
		.out_row (out_row_4_3),
		.out_col (out_col_4_3),
		.out_data (out_data_4_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_4;
	wire signed [DATA_WIDTH-1:0] out_col_4_4;
	wire signed [DATA_WIDTH-1:0] out_data_4_4;
	integer_mac_pe mac_pe_4_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_3),
		.in_col (out_col_3_4),
		.out_row (out_row_4_4),
		.out_col (out_col_4_4),
		.out_data (out_data_4_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_5;
	wire signed [DATA_WIDTH-1:0] out_col_4_5;
	wire signed [DATA_WIDTH-1:0] out_data_4_5;
	integer_mac_pe mac_pe_4_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_4),
		.in_col (out_col_3_5),
		.out_row (out_row_4_5),
		.out_col (out_col_4_5),
		.out_data (out_data_4_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_6;
	wire signed [DATA_WIDTH-1:0] out_col_4_6;
	wire signed [DATA_WIDTH-1:0] out_data_4_6;
	integer_mac_pe mac_pe_4_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_5),
		.in_col (out_col_3_6),
		.out_row (out_row_4_6),
		.out_col (out_col_4_6),
		.out_data (out_data_4_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_7;
	wire signed [DATA_WIDTH-1:0] out_col_4_7;
	wire signed [DATA_WIDTH-1:0] out_data_4_7;
	integer_mac_pe mac_pe_4_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_6),
		.in_col (out_col_3_7),
		.out_row (out_row_4_7),
		.out_col (out_col_4_7),
		.out_data (out_data_4_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_8;
	wire signed [DATA_WIDTH-1:0] out_col_4_8;
	wire signed [DATA_WIDTH-1:0] out_data_4_8;
	integer_mac_pe mac_pe_4_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_7),
		.in_col (out_col_3_8),
		.out_row (out_row_4_8),
		.out_col (out_col_4_8),
		.out_data (out_data_4_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_9;
	wire signed [DATA_WIDTH-1:0] out_col_4_9;
	wire signed [DATA_WIDTH-1:0] out_data_4_9;
	integer_mac_pe mac_pe_4_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_8),
		.in_col (out_col_3_9),
		.out_row (out_row_4_9),
		.out_col (out_col_4_9),
		.out_data (out_data_4_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_10;
	wire signed [DATA_WIDTH-1:0] out_col_4_10;
	wire signed [DATA_WIDTH-1:0] out_data_4_10;
	integer_mac_pe mac_pe_4_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_9),
		.in_col (out_col_3_10),
		.out_row (out_row_4_10),
		.out_col (out_col_4_10),
		.out_data (out_data_4_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_11;
	wire signed [DATA_WIDTH-1:0] out_col_4_11;
	wire signed [DATA_WIDTH-1:0] out_data_4_11;
	integer_mac_pe mac_pe_4_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_10),
		.in_col (out_col_3_11),
		.out_row (out_row_4_11),
		.out_col (out_col_4_11),
		.out_data (out_data_4_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_12;
	wire signed [DATA_WIDTH-1:0] out_col_4_12;
	wire signed [DATA_WIDTH-1:0] out_data_4_12;
	integer_mac_pe mac_pe_4_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_11),
		.in_col (out_col_3_12),
		.out_row (out_row_4_12),
		.out_col (out_col_4_12),
		.out_data (out_data_4_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_13;
	wire signed [DATA_WIDTH-1:0] out_col_4_13;
	wire signed [DATA_WIDTH-1:0] out_data_4_13;
	integer_mac_pe mac_pe_4_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_12),
		.in_col (out_col_3_13),
		.out_row (out_row_4_13),
		.out_col (out_col_4_13),
		.out_data (out_data_4_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_14;
	wire signed [DATA_WIDTH-1:0] out_col_4_14;
	wire signed [DATA_WIDTH-1:0] out_data_4_14;
	integer_mac_pe mac_pe_4_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_13),
		.in_col (out_col_3_14),
		.out_row (out_row_4_14),
		.out_col (out_col_4_14),
		.out_data (out_data_4_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_15;
	wire signed [DATA_WIDTH-1:0] out_col_4_15;
	wire signed [DATA_WIDTH-1:0] out_data_4_15;
	integer_mac_pe mac_pe_4_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_14),
		.in_col (out_col_3_15),
		.out_row (out_row_4_15),
		.out_col (out_col_4_15),
		.out_data (out_data_4_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_16;
	wire signed [DATA_WIDTH-1:0] out_col_4_16;
	wire signed [DATA_WIDTH-1:0] out_data_4_16;
	integer_mac_pe mac_pe_4_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_15),
		.in_col (out_col_3_16),
		.out_row (out_row_4_16),
		.out_col (out_col_4_16),
		.out_data (out_data_4_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_17;
	wire signed [DATA_WIDTH-1:0] out_col_4_17;
	wire signed [DATA_WIDTH-1:0] out_data_4_17;
	integer_mac_pe mac_pe_4_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_16),
		.in_col (out_col_3_17),
		.out_row (out_row_4_17),
		.out_col (out_col_4_17),
		.out_data (out_data_4_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_18;
	wire signed [DATA_WIDTH-1:0] out_col_4_18;
	wire signed [DATA_WIDTH-1:0] out_data_4_18;
	integer_mac_pe mac_pe_4_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_17),
		.in_col (out_col_3_18),
		.out_row (out_row_4_18),
		.out_col (out_col_4_18),
		.out_data (out_data_4_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_19;
	wire signed [DATA_WIDTH-1:0] out_col_4_19;
	wire signed [DATA_WIDTH-1:0] out_data_4_19;
	integer_mac_pe mac_pe_4_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_18),
		.in_col (out_col_3_19),
		.out_row (out_row_4_19),
		.out_col (out_col_4_19),
		.out_data (out_data_4_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_20;
	wire signed [DATA_WIDTH-1:0] out_col_4_20;
	wire signed [DATA_WIDTH-1:0] out_data_4_20;
	integer_mac_pe mac_pe_4_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_19),
		.in_col (out_col_3_20),
		.out_row (out_row_4_20),
		.out_col (out_col_4_20),
		.out_data (out_data_4_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_21;
	wire signed [DATA_WIDTH-1:0] out_col_4_21;
	wire signed [DATA_WIDTH-1:0] out_data_4_21;
	integer_mac_pe mac_pe_4_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_20),
		.in_col (out_col_3_21),
		.out_row (out_row_4_21),
		.out_col (out_col_4_21),
		.out_data (out_data_4_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_22;
	wire signed [DATA_WIDTH-1:0] out_col_4_22;
	wire signed [DATA_WIDTH-1:0] out_data_4_22;
	integer_mac_pe mac_pe_4_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_21),
		.in_col (out_col_3_22),
		.out_row (out_row_4_22),
		.out_col (out_col_4_22),
		.out_data (out_data_4_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_23;
	wire signed [DATA_WIDTH-1:0] out_col_4_23;
	wire signed [DATA_WIDTH-1:0] out_data_4_23;
	integer_mac_pe mac_pe_4_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_22),
		.in_col (out_col_3_23),
		.out_row (out_row_4_23),
		.out_col (out_col_4_23),
		.out_data (out_data_4_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_24;
	wire signed [DATA_WIDTH-1:0] out_col_4_24;
	wire signed [DATA_WIDTH-1:0] out_data_4_24;
	integer_mac_pe mac_pe_4_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_23),
		.in_col (out_col_3_24),
		.out_row (out_row_4_24),
		.out_col (out_col_4_24),
		.out_data (out_data_4_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_25;
	wire signed [DATA_WIDTH-1:0] out_col_4_25;
	wire signed [DATA_WIDTH-1:0] out_data_4_25;
	integer_mac_pe mac_pe_4_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_24),
		.in_col (out_col_3_25),
		.out_row (out_row_4_25),
		.out_col (out_col_4_25),
		.out_data (out_data_4_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_26;
	wire signed [DATA_WIDTH-1:0] out_col_4_26;
	wire signed [DATA_WIDTH-1:0] out_data_4_26;
	integer_mac_pe mac_pe_4_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_25),
		.in_col (out_col_3_26),
		.out_row (out_row_4_26),
		.out_col (out_col_4_26),
		.out_data (out_data_4_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_27;
	wire signed [DATA_WIDTH-1:0] out_col_4_27;
	wire signed [DATA_WIDTH-1:0] out_data_4_27;
	integer_mac_pe mac_pe_4_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_26),
		.in_col (out_col_3_27),
		.out_row (out_row_4_27),
		.out_col (out_col_4_27),
		.out_data (out_data_4_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_28;
	wire signed [DATA_WIDTH-1:0] out_col_4_28;
	wire signed [DATA_WIDTH-1:0] out_data_4_28;
	integer_mac_pe mac_pe_4_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_27),
		.in_col (out_col_3_28),
		.out_row (out_row_4_28),
		.out_col (out_col_4_28),
		.out_data (out_data_4_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_29;
	wire signed [DATA_WIDTH-1:0] out_col_4_29;
	wire signed [DATA_WIDTH-1:0] out_data_4_29;
	integer_mac_pe mac_pe_4_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_28),
		.in_col (out_col_3_29),
		.out_row (out_row_4_29),
		.out_col (out_col_4_29),
		.out_data (out_data_4_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_30;
	wire signed [DATA_WIDTH-1:0] out_col_4_30;
	wire signed [DATA_WIDTH-1:0] out_data_4_30;
	integer_mac_pe mac_pe_4_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_29),
		.in_col (out_col_3_30),
		.out_row (out_row_4_30),
		.out_col (out_col_4_30),
		.out_data (out_data_4_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_4_31;
	wire signed [DATA_WIDTH-1:0] out_col_4_31;
	wire signed [DATA_WIDTH-1:0] out_data_4_31;
	integer_mac_pe mac_pe_4_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_4_30),
		.in_col (out_col_3_31),
		.out_row (out_row_4_31),
		.out_col (out_col_4_31),
		.out_data (out_data_4_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_0;
	wire signed [DATA_WIDTH-1:0] out_col_5_0;
	wire signed [DATA_WIDTH-1:0] out_data_5_0;
	integer_mac_pe mac_pe_5_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_5_out),
		.in_col (out_col_4_0),
		.out_row (out_row_5_0),
		.out_col (out_col_5_0),
		.out_data (out_data_5_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_1;
	wire signed [DATA_WIDTH-1:0] out_col_5_1;
	wire signed [DATA_WIDTH-1:0] out_data_5_1;
	integer_mac_pe mac_pe_5_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_0),
		.in_col (out_col_4_1),
		.out_row (out_row_5_1),
		.out_col (out_col_5_1),
		.out_data (out_data_5_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_2;
	wire signed [DATA_WIDTH-1:0] out_col_5_2;
	wire signed [DATA_WIDTH-1:0] out_data_5_2;
	integer_mac_pe mac_pe_5_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_1),
		.in_col (out_col_4_2),
		.out_row (out_row_5_2),
		.out_col (out_col_5_2),
		.out_data (out_data_5_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_3;
	wire signed [DATA_WIDTH-1:0] out_col_5_3;
	wire signed [DATA_WIDTH-1:0] out_data_5_3;
	integer_mac_pe mac_pe_5_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_2),
		.in_col (out_col_4_3),
		.out_row (out_row_5_3),
		.out_col (out_col_5_3),
		.out_data (out_data_5_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_4;
	wire signed [DATA_WIDTH-1:0] out_col_5_4;
	wire signed [DATA_WIDTH-1:0] out_data_5_4;
	integer_mac_pe mac_pe_5_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_3),
		.in_col (out_col_4_4),
		.out_row (out_row_5_4),
		.out_col (out_col_5_4),
		.out_data (out_data_5_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_5;
	wire signed [DATA_WIDTH-1:0] out_col_5_5;
	wire signed [DATA_WIDTH-1:0] out_data_5_5;
	integer_mac_pe mac_pe_5_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_4),
		.in_col (out_col_4_5),
		.out_row (out_row_5_5),
		.out_col (out_col_5_5),
		.out_data (out_data_5_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_6;
	wire signed [DATA_WIDTH-1:0] out_col_5_6;
	wire signed [DATA_WIDTH-1:0] out_data_5_6;
	integer_mac_pe mac_pe_5_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_5),
		.in_col (out_col_4_6),
		.out_row (out_row_5_6),
		.out_col (out_col_5_6),
		.out_data (out_data_5_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_7;
	wire signed [DATA_WIDTH-1:0] out_col_5_7;
	wire signed [DATA_WIDTH-1:0] out_data_5_7;
	integer_mac_pe mac_pe_5_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_6),
		.in_col (out_col_4_7),
		.out_row (out_row_5_7),
		.out_col (out_col_5_7),
		.out_data (out_data_5_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_8;
	wire signed [DATA_WIDTH-1:0] out_col_5_8;
	wire signed [DATA_WIDTH-1:0] out_data_5_8;
	integer_mac_pe mac_pe_5_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_7),
		.in_col (out_col_4_8),
		.out_row (out_row_5_8),
		.out_col (out_col_5_8),
		.out_data (out_data_5_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_9;
	wire signed [DATA_WIDTH-1:0] out_col_5_9;
	wire signed [DATA_WIDTH-1:0] out_data_5_9;
	integer_mac_pe mac_pe_5_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_8),
		.in_col (out_col_4_9),
		.out_row (out_row_5_9),
		.out_col (out_col_5_9),
		.out_data (out_data_5_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_10;
	wire signed [DATA_WIDTH-1:0] out_col_5_10;
	wire signed [DATA_WIDTH-1:0] out_data_5_10;
	integer_mac_pe mac_pe_5_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_9),
		.in_col (out_col_4_10),
		.out_row (out_row_5_10),
		.out_col (out_col_5_10),
		.out_data (out_data_5_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_11;
	wire signed [DATA_WIDTH-1:0] out_col_5_11;
	wire signed [DATA_WIDTH-1:0] out_data_5_11;
	integer_mac_pe mac_pe_5_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_10),
		.in_col (out_col_4_11),
		.out_row (out_row_5_11),
		.out_col (out_col_5_11),
		.out_data (out_data_5_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_12;
	wire signed [DATA_WIDTH-1:0] out_col_5_12;
	wire signed [DATA_WIDTH-1:0] out_data_5_12;
	integer_mac_pe mac_pe_5_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_11),
		.in_col (out_col_4_12),
		.out_row (out_row_5_12),
		.out_col (out_col_5_12),
		.out_data (out_data_5_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_13;
	wire signed [DATA_WIDTH-1:0] out_col_5_13;
	wire signed [DATA_WIDTH-1:0] out_data_5_13;
	integer_mac_pe mac_pe_5_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_12),
		.in_col (out_col_4_13),
		.out_row (out_row_5_13),
		.out_col (out_col_5_13),
		.out_data (out_data_5_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_14;
	wire signed [DATA_WIDTH-1:0] out_col_5_14;
	wire signed [DATA_WIDTH-1:0] out_data_5_14;
	integer_mac_pe mac_pe_5_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_13),
		.in_col (out_col_4_14),
		.out_row (out_row_5_14),
		.out_col (out_col_5_14),
		.out_data (out_data_5_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_15;
	wire signed [DATA_WIDTH-1:0] out_col_5_15;
	wire signed [DATA_WIDTH-1:0] out_data_5_15;
	integer_mac_pe mac_pe_5_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_14),
		.in_col (out_col_4_15),
		.out_row (out_row_5_15),
		.out_col (out_col_5_15),
		.out_data (out_data_5_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_16;
	wire signed [DATA_WIDTH-1:0] out_col_5_16;
	wire signed [DATA_WIDTH-1:0] out_data_5_16;
	integer_mac_pe mac_pe_5_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_15),
		.in_col (out_col_4_16),
		.out_row (out_row_5_16),
		.out_col (out_col_5_16),
		.out_data (out_data_5_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_17;
	wire signed [DATA_WIDTH-1:0] out_col_5_17;
	wire signed [DATA_WIDTH-1:0] out_data_5_17;
	integer_mac_pe mac_pe_5_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_16),
		.in_col (out_col_4_17),
		.out_row (out_row_5_17),
		.out_col (out_col_5_17),
		.out_data (out_data_5_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_18;
	wire signed [DATA_WIDTH-1:0] out_col_5_18;
	wire signed [DATA_WIDTH-1:0] out_data_5_18;
	integer_mac_pe mac_pe_5_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_17),
		.in_col (out_col_4_18),
		.out_row (out_row_5_18),
		.out_col (out_col_5_18),
		.out_data (out_data_5_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_19;
	wire signed [DATA_WIDTH-1:0] out_col_5_19;
	wire signed [DATA_WIDTH-1:0] out_data_5_19;
	integer_mac_pe mac_pe_5_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_18),
		.in_col (out_col_4_19),
		.out_row (out_row_5_19),
		.out_col (out_col_5_19),
		.out_data (out_data_5_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_20;
	wire signed [DATA_WIDTH-1:0] out_col_5_20;
	wire signed [DATA_WIDTH-1:0] out_data_5_20;
	integer_mac_pe mac_pe_5_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_19),
		.in_col (out_col_4_20),
		.out_row (out_row_5_20),
		.out_col (out_col_5_20),
		.out_data (out_data_5_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_21;
	wire signed [DATA_WIDTH-1:0] out_col_5_21;
	wire signed [DATA_WIDTH-1:0] out_data_5_21;
	integer_mac_pe mac_pe_5_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_20),
		.in_col (out_col_4_21),
		.out_row (out_row_5_21),
		.out_col (out_col_5_21),
		.out_data (out_data_5_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_22;
	wire signed [DATA_WIDTH-1:0] out_col_5_22;
	wire signed [DATA_WIDTH-1:0] out_data_5_22;
	integer_mac_pe mac_pe_5_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_21),
		.in_col (out_col_4_22),
		.out_row (out_row_5_22),
		.out_col (out_col_5_22),
		.out_data (out_data_5_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_23;
	wire signed [DATA_WIDTH-1:0] out_col_5_23;
	wire signed [DATA_WIDTH-1:0] out_data_5_23;
	integer_mac_pe mac_pe_5_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_22),
		.in_col (out_col_4_23),
		.out_row (out_row_5_23),
		.out_col (out_col_5_23),
		.out_data (out_data_5_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_24;
	wire signed [DATA_WIDTH-1:0] out_col_5_24;
	wire signed [DATA_WIDTH-1:0] out_data_5_24;
	integer_mac_pe mac_pe_5_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_23),
		.in_col (out_col_4_24),
		.out_row (out_row_5_24),
		.out_col (out_col_5_24),
		.out_data (out_data_5_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_25;
	wire signed [DATA_WIDTH-1:0] out_col_5_25;
	wire signed [DATA_WIDTH-1:0] out_data_5_25;
	integer_mac_pe mac_pe_5_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_24),
		.in_col (out_col_4_25),
		.out_row (out_row_5_25),
		.out_col (out_col_5_25),
		.out_data (out_data_5_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_26;
	wire signed [DATA_WIDTH-1:0] out_col_5_26;
	wire signed [DATA_WIDTH-1:0] out_data_5_26;
	integer_mac_pe mac_pe_5_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_25),
		.in_col (out_col_4_26),
		.out_row (out_row_5_26),
		.out_col (out_col_5_26),
		.out_data (out_data_5_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_27;
	wire signed [DATA_WIDTH-1:0] out_col_5_27;
	wire signed [DATA_WIDTH-1:0] out_data_5_27;
	integer_mac_pe mac_pe_5_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_26),
		.in_col (out_col_4_27),
		.out_row (out_row_5_27),
		.out_col (out_col_5_27),
		.out_data (out_data_5_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_28;
	wire signed [DATA_WIDTH-1:0] out_col_5_28;
	wire signed [DATA_WIDTH-1:0] out_data_5_28;
	integer_mac_pe mac_pe_5_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_27),
		.in_col (out_col_4_28),
		.out_row (out_row_5_28),
		.out_col (out_col_5_28),
		.out_data (out_data_5_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_29;
	wire signed [DATA_WIDTH-1:0] out_col_5_29;
	wire signed [DATA_WIDTH-1:0] out_data_5_29;
	integer_mac_pe mac_pe_5_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_28),
		.in_col (out_col_4_29),
		.out_row (out_row_5_29),
		.out_col (out_col_5_29),
		.out_data (out_data_5_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_30;
	wire signed [DATA_WIDTH-1:0] out_col_5_30;
	wire signed [DATA_WIDTH-1:0] out_data_5_30;
	integer_mac_pe mac_pe_5_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_29),
		.in_col (out_col_4_30),
		.out_row (out_row_5_30),
		.out_col (out_col_5_30),
		.out_data (out_data_5_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_5_31;
	wire signed [DATA_WIDTH-1:0] out_col_5_31;
	wire signed [DATA_WIDTH-1:0] out_data_5_31;
	integer_mac_pe mac_pe_5_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_5_30),
		.in_col (out_col_4_31),
		.out_row (out_row_5_31),
		.out_col (out_col_5_31),
		.out_data (out_data_5_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_0;
	wire signed [DATA_WIDTH-1:0] out_col_6_0;
	wire signed [DATA_WIDTH-1:0] out_data_6_0;
	integer_mac_pe mac_pe_6_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_6_out),
		.in_col (out_col_5_0),
		.out_row (out_row_6_0),
		.out_col (out_col_6_0),
		.out_data (out_data_6_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_1;
	wire signed [DATA_WIDTH-1:0] out_col_6_1;
	wire signed [DATA_WIDTH-1:0] out_data_6_1;
	integer_mac_pe mac_pe_6_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_0),
		.in_col (out_col_5_1),
		.out_row (out_row_6_1),
		.out_col (out_col_6_1),
		.out_data (out_data_6_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_2;
	wire signed [DATA_WIDTH-1:0] out_col_6_2;
	wire signed [DATA_WIDTH-1:0] out_data_6_2;
	integer_mac_pe mac_pe_6_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_1),
		.in_col (out_col_5_2),
		.out_row (out_row_6_2),
		.out_col (out_col_6_2),
		.out_data (out_data_6_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_3;
	wire signed [DATA_WIDTH-1:0] out_col_6_3;
	wire signed [DATA_WIDTH-1:0] out_data_6_3;
	integer_mac_pe mac_pe_6_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_2),
		.in_col (out_col_5_3),
		.out_row (out_row_6_3),
		.out_col (out_col_6_3),
		.out_data (out_data_6_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_4;
	wire signed [DATA_WIDTH-1:0] out_col_6_4;
	wire signed [DATA_WIDTH-1:0] out_data_6_4;
	integer_mac_pe mac_pe_6_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_3),
		.in_col (out_col_5_4),
		.out_row (out_row_6_4),
		.out_col (out_col_6_4),
		.out_data (out_data_6_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_5;
	wire signed [DATA_WIDTH-1:0] out_col_6_5;
	wire signed [DATA_WIDTH-1:0] out_data_6_5;
	integer_mac_pe mac_pe_6_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_4),
		.in_col (out_col_5_5),
		.out_row (out_row_6_5),
		.out_col (out_col_6_5),
		.out_data (out_data_6_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_6;
	wire signed [DATA_WIDTH-1:0] out_col_6_6;
	wire signed [DATA_WIDTH-1:0] out_data_6_6;
	integer_mac_pe mac_pe_6_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_5),
		.in_col (out_col_5_6),
		.out_row (out_row_6_6),
		.out_col (out_col_6_6),
		.out_data (out_data_6_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_7;
	wire signed [DATA_WIDTH-1:0] out_col_6_7;
	wire signed [DATA_WIDTH-1:0] out_data_6_7;
	integer_mac_pe mac_pe_6_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_6),
		.in_col (out_col_5_7),
		.out_row (out_row_6_7),
		.out_col (out_col_6_7),
		.out_data (out_data_6_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_8;
	wire signed [DATA_WIDTH-1:0] out_col_6_8;
	wire signed [DATA_WIDTH-1:0] out_data_6_8;
	integer_mac_pe mac_pe_6_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_7),
		.in_col (out_col_5_8),
		.out_row (out_row_6_8),
		.out_col (out_col_6_8),
		.out_data (out_data_6_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_9;
	wire signed [DATA_WIDTH-1:0] out_col_6_9;
	wire signed [DATA_WIDTH-1:0] out_data_6_9;
	integer_mac_pe mac_pe_6_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_8),
		.in_col (out_col_5_9),
		.out_row (out_row_6_9),
		.out_col (out_col_6_9),
		.out_data (out_data_6_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_10;
	wire signed [DATA_WIDTH-1:0] out_col_6_10;
	wire signed [DATA_WIDTH-1:0] out_data_6_10;
	integer_mac_pe mac_pe_6_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_9),
		.in_col (out_col_5_10),
		.out_row (out_row_6_10),
		.out_col (out_col_6_10),
		.out_data (out_data_6_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_11;
	wire signed [DATA_WIDTH-1:0] out_col_6_11;
	wire signed [DATA_WIDTH-1:0] out_data_6_11;
	integer_mac_pe mac_pe_6_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_10),
		.in_col (out_col_5_11),
		.out_row (out_row_6_11),
		.out_col (out_col_6_11),
		.out_data (out_data_6_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_12;
	wire signed [DATA_WIDTH-1:0] out_col_6_12;
	wire signed [DATA_WIDTH-1:0] out_data_6_12;
	integer_mac_pe mac_pe_6_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_11),
		.in_col (out_col_5_12),
		.out_row (out_row_6_12),
		.out_col (out_col_6_12),
		.out_data (out_data_6_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_13;
	wire signed [DATA_WIDTH-1:0] out_col_6_13;
	wire signed [DATA_WIDTH-1:0] out_data_6_13;
	integer_mac_pe mac_pe_6_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_12),
		.in_col (out_col_5_13),
		.out_row (out_row_6_13),
		.out_col (out_col_6_13),
		.out_data (out_data_6_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_14;
	wire signed [DATA_WIDTH-1:0] out_col_6_14;
	wire signed [DATA_WIDTH-1:0] out_data_6_14;
	integer_mac_pe mac_pe_6_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_13),
		.in_col (out_col_5_14),
		.out_row (out_row_6_14),
		.out_col (out_col_6_14),
		.out_data (out_data_6_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_15;
	wire signed [DATA_WIDTH-1:0] out_col_6_15;
	wire signed [DATA_WIDTH-1:0] out_data_6_15;
	integer_mac_pe mac_pe_6_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_14),
		.in_col (out_col_5_15),
		.out_row (out_row_6_15),
		.out_col (out_col_6_15),
		.out_data (out_data_6_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_16;
	wire signed [DATA_WIDTH-1:0] out_col_6_16;
	wire signed [DATA_WIDTH-1:0] out_data_6_16;
	integer_mac_pe mac_pe_6_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_15),
		.in_col (out_col_5_16),
		.out_row (out_row_6_16),
		.out_col (out_col_6_16),
		.out_data (out_data_6_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_17;
	wire signed [DATA_WIDTH-1:0] out_col_6_17;
	wire signed [DATA_WIDTH-1:0] out_data_6_17;
	integer_mac_pe mac_pe_6_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_16),
		.in_col (out_col_5_17),
		.out_row (out_row_6_17),
		.out_col (out_col_6_17),
		.out_data (out_data_6_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_18;
	wire signed [DATA_WIDTH-1:0] out_col_6_18;
	wire signed [DATA_WIDTH-1:0] out_data_6_18;
	integer_mac_pe mac_pe_6_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_17),
		.in_col (out_col_5_18),
		.out_row (out_row_6_18),
		.out_col (out_col_6_18),
		.out_data (out_data_6_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_19;
	wire signed [DATA_WIDTH-1:0] out_col_6_19;
	wire signed [DATA_WIDTH-1:0] out_data_6_19;
	integer_mac_pe mac_pe_6_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_18),
		.in_col (out_col_5_19),
		.out_row (out_row_6_19),
		.out_col (out_col_6_19),
		.out_data (out_data_6_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_20;
	wire signed [DATA_WIDTH-1:0] out_col_6_20;
	wire signed [DATA_WIDTH-1:0] out_data_6_20;
	integer_mac_pe mac_pe_6_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_19),
		.in_col (out_col_5_20),
		.out_row (out_row_6_20),
		.out_col (out_col_6_20),
		.out_data (out_data_6_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_21;
	wire signed [DATA_WIDTH-1:0] out_col_6_21;
	wire signed [DATA_WIDTH-1:0] out_data_6_21;
	integer_mac_pe mac_pe_6_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_20),
		.in_col (out_col_5_21),
		.out_row (out_row_6_21),
		.out_col (out_col_6_21),
		.out_data (out_data_6_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_22;
	wire signed [DATA_WIDTH-1:0] out_col_6_22;
	wire signed [DATA_WIDTH-1:0] out_data_6_22;
	integer_mac_pe mac_pe_6_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_21),
		.in_col (out_col_5_22),
		.out_row (out_row_6_22),
		.out_col (out_col_6_22),
		.out_data (out_data_6_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_23;
	wire signed [DATA_WIDTH-1:0] out_col_6_23;
	wire signed [DATA_WIDTH-1:0] out_data_6_23;
	integer_mac_pe mac_pe_6_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_22),
		.in_col (out_col_5_23),
		.out_row (out_row_6_23),
		.out_col (out_col_6_23),
		.out_data (out_data_6_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_24;
	wire signed [DATA_WIDTH-1:0] out_col_6_24;
	wire signed [DATA_WIDTH-1:0] out_data_6_24;
	integer_mac_pe mac_pe_6_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_23),
		.in_col (out_col_5_24),
		.out_row (out_row_6_24),
		.out_col (out_col_6_24),
		.out_data (out_data_6_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_25;
	wire signed [DATA_WIDTH-1:0] out_col_6_25;
	wire signed [DATA_WIDTH-1:0] out_data_6_25;
	integer_mac_pe mac_pe_6_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_24),
		.in_col (out_col_5_25),
		.out_row (out_row_6_25),
		.out_col (out_col_6_25),
		.out_data (out_data_6_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_26;
	wire signed [DATA_WIDTH-1:0] out_col_6_26;
	wire signed [DATA_WIDTH-1:0] out_data_6_26;
	integer_mac_pe mac_pe_6_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_25),
		.in_col (out_col_5_26),
		.out_row (out_row_6_26),
		.out_col (out_col_6_26),
		.out_data (out_data_6_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_27;
	wire signed [DATA_WIDTH-1:0] out_col_6_27;
	wire signed [DATA_WIDTH-1:0] out_data_6_27;
	integer_mac_pe mac_pe_6_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_26),
		.in_col (out_col_5_27),
		.out_row (out_row_6_27),
		.out_col (out_col_6_27),
		.out_data (out_data_6_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_28;
	wire signed [DATA_WIDTH-1:0] out_col_6_28;
	wire signed [DATA_WIDTH-1:0] out_data_6_28;
	integer_mac_pe mac_pe_6_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_27),
		.in_col (out_col_5_28),
		.out_row (out_row_6_28),
		.out_col (out_col_6_28),
		.out_data (out_data_6_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_29;
	wire signed [DATA_WIDTH-1:0] out_col_6_29;
	wire signed [DATA_WIDTH-1:0] out_data_6_29;
	integer_mac_pe mac_pe_6_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_28),
		.in_col (out_col_5_29),
		.out_row (out_row_6_29),
		.out_col (out_col_6_29),
		.out_data (out_data_6_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_30;
	wire signed [DATA_WIDTH-1:0] out_col_6_30;
	wire signed [DATA_WIDTH-1:0] out_data_6_30;
	integer_mac_pe mac_pe_6_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_29),
		.in_col (out_col_5_30),
		.out_row (out_row_6_30),
		.out_col (out_col_6_30),
		.out_data (out_data_6_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_6_31;
	wire signed [DATA_WIDTH-1:0] out_col_6_31;
	wire signed [DATA_WIDTH-1:0] out_data_6_31;
	integer_mac_pe mac_pe_6_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_6_30),
		.in_col (out_col_5_31),
		.out_row (out_row_6_31),
		.out_col (out_col_6_31),
		.out_data (out_data_6_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_0;
	wire signed [DATA_WIDTH-1:0] out_col_7_0;
	wire signed [DATA_WIDTH-1:0] out_data_7_0;
	integer_mac_pe mac_pe_7_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_7_out),
		.in_col (out_col_6_0),
		.out_row (out_row_7_0),
		.out_col (out_col_7_0),
		.out_data (out_data_7_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_1;
	wire signed [DATA_WIDTH-1:0] out_col_7_1;
	wire signed [DATA_WIDTH-1:0] out_data_7_1;
	integer_mac_pe mac_pe_7_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_0),
		.in_col (out_col_6_1),
		.out_row (out_row_7_1),
		.out_col (out_col_7_1),
		.out_data (out_data_7_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_2;
	wire signed [DATA_WIDTH-1:0] out_col_7_2;
	wire signed [DATA_WIDTH-1:0] out_data_7_2;
	integer_mac_pe mac_pe_7_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_1),
		.in_col (out_col_6_2),
		.out_row (out_row_7_2),
		.out_col (out_col_7_2),
		.out_data (out_data_7_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_3;
	wire signed [DATA_WIDTH-1:0] out_col_7_3;
	wire signed [DATA_WIDTH-1:0] out_data_7_3;
	integer_mac_pe mac_pe_7_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_2),
		.in_col (out_col_6_3),
		.out_row (out_row_7_3),
		.out_col (out_col_7_3),
		.out_data (out_data_7_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_4;
	wire signed [DATA_WIDTH-1:0] out_col_7_4;
	wire signed [DATA_WIDTH-1:0] out_data_7_4;
	integer_mac_pe mac_pe_7_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_3),
		.in_col (out_col_6_4),
		.out_row (out_row_7_4),
		.out_col (out_col_7_4),
		.out_data (out_data_7_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_5;
	wire signed [DATA_WIDTH-1:0] out_col_7_5;
	wire signed [DATA_WIDTH-1:0] out_data_7_5;
	integer_mac_pe mac_pe_7_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_4),
		.in_col (out_col_6_5),
		.out_row (out_row_7_5),
		.out_col (out_col_7_5),
		.out_data (out_data_7_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_6;
	wire signed [DATA_WIDTH-1:0] out_col_7_6;
	wire signed [DATA_WIDTH-1:0] out_data_7_6;
	integer_mac_pe mac_pe_7_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_5),
		.in_col (out_col_6_6),
		.out_row (out_row_7_6),
		.out_col (out_col_7_6),
		.out_data (out_data_7_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_7;
	wire signed [DATA_WIDTH-1:0] out_col_7_7;
	wire signed [DATA_WIDTH-1:0] out_data_7_7;
	integer_mac_pe mac_pe_7_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_6),
		.in_col (out_col_6_7),
		.out_row (out_row_7_7),
		.out_col (out_col_7_7),
		.out_data (out_data_7_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_8;
	wire signed [DATA_WIDTH-1:0] out_col_7_8;
	wire signed [DATA_WIDTH-1:0] out_data_7_8;
	integer_mac_pe mac_pe_7_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_7),
		.in_col (out_col_6_8),
		.out_row (out_row_7_8),
		.out_col (out_col_7_8),
		.out_data (out_data_7_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_9;
	wire signed [DATA_WIDTH-1:0] out_col_7_9;
	wire signed [DATA_WIDTH-1:0] out_data_7_9;
	integer_mac_pe mac_pe_7_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_8),
		.in_col (out_col_6_9),
		.out_row (out_row_7_9),
		.out_col (out_col_7_9),
		.out_data (out_data_7_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_10;
	wire signed [DATA_WIDTH-1:0] out_col_7_10;
	wire signed [DATA_WIDTH-1:0] out_data_7_10;
	integer_mac_pe mac_pe_7_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_9),
		.in_col (out_col_6_10),
		.out_row (out_row_7_10),
		.out_col (out_col_7_10),
		.out_data (out_data_7_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_11;
	wire signed [DATA_WIDTH-1:0] out_col_7_11;
	wire signed [DATA_WIDTH-1:0] out_data_7_11;
	integer_mac_pe mac_pe_7_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_10),
		.in_col (out_col_6_11),
		.out_row (out_row_7_11),
		.out_col (out_col_7_11),
		.out_data (out_data_7_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_12;
	wire signed [DATA_WIDTH-1:0] out_col_7_12;
	wire signed [DATA_WIDTH-1:0] out_data_7_12;
	integer_mac_pe mac_pe_7_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_11),
		.in_col (out_col_6_12),
		.out_row (out_row_7_12),
		.out_col (out_col_7_12),
		.out_data (out_data_7_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_13;
	wire signed [DATA_WIDTH-1:0] out_col_7_13;
	wire signed [DATA_WIDTH-1:0] out_data_7_13;
	integer_mac_pe mac_pe_7_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_12),
		.in_col (out_col_6_13),
		.out_row (out_row_7_13),
		.out_col (out_col_7_13),
		.out_data (out_data_7_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_14;
	wire signed [DATA_WIDTH-1:0] out_col_7_14;
	wire signed [DATA_WIDTH-1:0] out_data_7_14;
	integer_mac_pe mac_pe_7_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_13),
		.in_col (out_col_6_14),
		.out_row (out_row_7_14),
		.out_col (out_col_7_14),
		.out_data (out_data_7_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_15;
	wire signed [DATA_WIDTH-1:0] out_col_7_15;
	wire signed [DATA_WIDTH-1:0] out_data_7_15;
	integer_mac_pe mac_pe_7_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_14),
		.in_col (out_col_6_15),
		.out_row (out_row_7_15),
		.out_col (out_col_7_15),
		.out_data (out_data_7_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_16;
	wire signed [DATA_WIDTH-1:0] out_col_7_16;
	wire signed [DATA_WIDTH-1:0] out_data_7_16;
	integer_mac_pe mac_pe_7_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_15),
		.in_col (out_col_6_16),
		.out_row (out_row_7_16),
		.out_col (out_col_7_16),
		.out_data (out_data_7_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_17;
	wire signed [DATA_WIDTH-1:0] out_col_7_17;
	wire signed [DATA_WIDTH-1:0] out_data_7_17;
	integer_mac_pe mac_pe_7_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_16),
		.in_col (out_col_6_17),
		.out_row (out_row_7_17),
		.out_col (out_col_7_17),
		.out_data (out_data_7_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_18;
	wire signed [DATA_WIDTH-1:0] out_col_7_18;
	wire signed [DATA_WIDTH-1:0] out_data_7_18;
	integer_mac_pe mac_pe_7_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_17),
		.in_col (out_col_6_18),
		.out_row (out_row_7_18),
		.out_col (out_col_7_18),
		.out_data (out_data_7_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_19;
	wire signed [DATA_WIDTH-1:0] out_col_7_19;
	wire signed [DATA_WIDTH-1:0] out_data_7_19;
	integer_mac_pe mac_pe_7_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_18),
		.in_col (out_col_6_19),
		.out_row (out_row_7_19),
		.out_col (out_col_7_19),
		.out_data (out_data_7_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_20;
	wire signed [DATA_WIDTH-1:0] out_col_7_20;
	wire signed [DATA_WIDTH-1:0] out_data_7_20;
	integer_mac_pe mac_pe_7_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_19),
		.in_col (out_col_6_20),
		.out_row (out_row_7_20),
		.out_col (out_col_7_20),
		.out_data (out_data_7_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_21;
	wire signed [DATA_WIDTH-1:0] out_col_7_21;
	wire signed [DATA_WIDTH-1:0] out_data_7_21;
	integer_mac_pe mac_pe_7_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_20),
		.in_col (out_col_6_21),
		.out_row (out_row_7_21),
		.out_col (out_col_7_21),
		.out_data (out_data_7_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_22;
	wire signed [DATA_WIDTH-1:0] out_col_7_22;
	wire signed [DATA_WIDTH-1:0] out_data_7_22;
	integer_mac_pe mac_pe_7_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_21),
		.in_col (out_col_6_22),
		.out_row (out_row_7_22),
		.out_col (out_col_7_22),
		.out_data (out_data_7_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_23;
	wire signed [DATA_WIDTH-1:0] out_col_7_23;
	wire signed [DATA_WIDTH-1:0] out_data_7_23;
	integer_mac_pe mac_pe_7_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_22),
		.in_col (out_col_6_23),
		.out_row (out_row_7_23),
		.out_col (out_col_7_23),
		.out_data (out_data_7_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_24;
	wire signed [DATA_WIDTH-1:0] out_col_7_24;
	wire signed [DATA_WIDTH-1:0] out_data_7_24;
	integer_mac_pe mac_pe_7_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_23),
		.in_col (out_col_6_24),
		.out_row (out_row_7_24),
		.out_col (out_col_7_24),
		.out_data (out_data_7_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_25;
	wire signed [DATA_WIDTH-1:0] out_col_7_25;
	wire signed [DATA_WIDTH-1:0] out_data_7_25;
	integer_mac_pe mac_pe_7_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_24),
		.in_col (out_col_6_25),
		.out_row (out_row_7_25),
		.out_col (out_col_7_25),
		.out_data (out_data_7_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_26;
	wire signed [DATA_WIDTH-1:0] out_col_7_26;
	wire signed [DATA_WIDTH-1:0] out_data_7_26;
	integer_mac_pe mac_pe_7_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_25),
		.in_col (out_col_6_26),
		.out_row (out_row_7_26),
		.out_col (out_col_7_26),
		.out_data (out_data_7_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_27;
	wire signed [DATA_WIDTH-1:0] out_col_7_27;
	wire signed [DATA_WIDTH-1:0] out_data_7_27;
	integer_mac_pe mac_pe_7_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_26),
		.in_col (out_col_6_27),
		.out_row (out_row_7_27),
		.out_col (out_col_7_27),
		.out_data (out_data_7_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_28;
	wire signed [DATA_WIDTH-1:0] out_col_7_28;
	wire signed [DATA_WIDTH-1:0] out_data_7_28;
	integer_mac_pe mac_pe_7_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_27),
		.in_col (out_col_6_28),
		.out_row (out_row_7_28),
		.out_col (out_col_7_28),
		.out_data (out_data_7_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_29;
	wire signed [DATA_WIDTH-1:0] out_col_7_29;
	wire signed [DATA_WIDTH-1:0] out_data_7_29;
	integer_mac_pe mac_pe_7_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_28),
		.in_col (out_col_6_29),
		.out_row (out_row_7_29),
		.out_col (out_col_7_29),
		.out_data (out_data_7_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_30;
	wire signed [DATA_WIDTH-1:0] out_col_7_30;
	wire signed [DATA_WIDTH-1:0] out_data_7_30;
	integer_mac_pe mac_pe_7_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_29),
		.in_col (out_col_6_30),
		.out_row (out_row_7_30),
		.out_col (out_col_7_30),
		.out_data (out_data_7_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_7_31;
	wire signed [DATA_WIDTH-1:0] out_col_7_31;
	wire signed [DATA_WIDTH-1:0] out_data_7_31;
	integer_mac_pe mac_pe_7_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_7_30),
		.in_col (out_col_6_31),
		.out_row (out_row_7_31),
		.out_col (out_col_7_31),
		.out_data (out_data_7_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_0;
	wire signed [DATA_WIDTH-1:0] out_col_8_0;
	wire signed [DATA_WIDTH-1:0] out_data_8_0;
	integer_mac_pe mac_pe_8_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_8_out),
		.in_col (out_col_7_0),
		.out_row (out_row_8_0),
		.out_col (out_col_8_0),
		.out_data (out_data_8_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_1;
	wire signed [DATA_WIDTH-1:0] out_col_8_1;
	wire signed [DATA_WIDTH-1:0] out_data_8_1;
	integer_mac_pe mac_pe_8_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_0),
		.in_col (out_col_7_1),
		.out_row (out_row_8_1),
		.out_col (out_col_8_1),
		.out_data (out_data_8_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_2;
	wire signed [DATA_WIDTH-1:0] out_col_8_2;
	wire signed [DATA_WIDTH-1:0] out_data_8_2;
	integer_mac_pe mac_pe_8_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_1),
		.in_col (out_col_7_2),
		.out_row (out_row_8_2),
		.out_col (out_col_8_2),
		.out_data (out_data_8_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_3;
	wire signed [DATA_WIDTH-1:0] out_col_8_3;
	wire signed [DATA_WIDTH-1:0] out_data_8_3;
	integer_mac_pe mac_pe_8_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_2),
		.in_col (out_col_7_3),
		.out_row (out_row_8_3),
		.out_col (out_col_8_3),
		.out_data (out_data_8_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_4;
	wire signed [DATA_WIDTH-1:0] out_col_8_4;
	wire signed [DATA_WIDTH-1:0] out_data_8_4;
	integer_mac_pe mac_pe_8_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_3),
		.in_col (out_col_7_4),
		.out_row (out_row_8_4),
		.out_col (out_col_8_4),
		.out_data (out_data_8_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_5;
	wire signed [DATA_WIDTH-1:0] out_col_8_5;
	wire signed [DATA_WIDTH-1:0] out_data_8_5;
	integer_mac_pe mac_pe_8_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_4),
		.in_col (out_col_7_5),
		.out_row (out_row_8_5),
		.out_col (out_col_8_5),
		.out_data (out_data_8_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_6;
	wire signed [DATA_WIDTH-1:0] out_col_8_6;
	wire signed [DATA_WIDTH-1:0] out_data_8_6;
	integer_mac_pe mac_pe_8_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_5),
		.in_col (out_col_7_6),
		.out_row (out_row_8_6),
		.out_col (out_col_8_6),
		.out_data (out_data_8_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_7;
	wire signed [DATA_WIDTH-1:0] out_col_8_7;
	wire signed [DATA_WIDTH-1:0] out_data_8_7;
	integer_mac_pe mac_pe_8_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_6),
		.in_col (out_col_7_7),
		.out_row (out_row_8_7),
		.out_col (out_col_8_7),
		.out_data (out_data_8_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_8;
	wire signed [DATA_WIDTH-1:0] out_col_8_8;
	wire signed [DATA_WIDTH-1:0] out_data_8_8;
	integer_mac_pe mac_pe_8_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_7),
		.in_col (out_col_7_8),
		.out_row (out_row_8_8),
		.out_col (out_col_8_8),
		.out_data (out_data_8_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_9;
	wire signed [DATA_WIDTH-1:0] out_col_8_9;
	wire signed [DATA_WIDTH-1:0] out_data_8_9;
	integer_mac_pe mac_pe_8_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_8),
		.in_col (out_col_7_9),
		.out_row (out_row_8_9),
		.out_col (out_col_8_9),
		.out_data (out_data_8_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_10;
	wire signed [DATA_WIDTH-1:0] out_col_8_10;
	wire signed [DATA_WIDTH-1:0] out_data_8_10;
	integer_mac_pe mac_pe_8_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_9),
		.in_col (out_col_7_10),
		.out_row (out_row_8_10),
		.out_col (out_col_8_10),
		.out_data (out_data_8_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_11;
	wire signed [DATA_WIDTH-1:0] out_col_8_11;
	wire signed [DATA_WIDTH-1:0] out_data_8_11;
	integer_mac_pe mac_pe_8_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_10),
		.in_col (out_col_7_11),
		.out_row (out_row_8_11),
		.out_col (out_col_8_11),
		.out_data (out_data_8_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_12;
	wire signed [DATA_WIDTH-1:0] out_col_8_12;
	wire signed [DATA_WIDTH-1:0] out_data_8_12;
	integer_mac_pe mac_pe_8_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_11),
		.in_col (out_col_7_12),
		.out_row (out_row_8_12),
		.out_col (out_col_8_12),
		.out_data (out_data_8_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_13;
	wire signed [DATA_WIDTH-1:0] out_col_8_13;
	wire signed [DATA_WIDTH-1:0] out_data_8_13;
	integer_mac_pe mac_pe_8_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_12),
		.in_col (out_col_7_13),
		.out_row (out_row_8_13),
		.out_col (out_col_8_13),
		.out_data (out_data_8_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_14;
	wire signed [DATA_WIDTH-1:0] out_col_8_14;
	wire signed [DATA_WIDTH-1:0] out_data_8_14;
	integer_mac_pe mac_pe_8_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_13),
		.in_col (out_col_7_14),
		.out_row (out_row_8_14),
		.out_col (out_col_8_14),
		.out_data (out_data_8_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_15;
	wire signed [DATA_WIDTH-1:0] out_col_8_15;
	wire signed [DATA_WIDTH-1:0] out_data_8_15;
	integer_mac_pe mac_pe_8_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_14),
		.in_col (out_col_7_15),
		.out_row (out_row_8_15),
		.out_col (out_col_8_15),
		.out_data (out_data_8_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_16;
	wire signed [DATA_WIDTH-1:0] out_col_8_16;
	wire signed [DATA_WIDTH-1:0] out_data_8_16;
	integer_mac_pe mac_pe_8_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_15),
		.in_col (out_col_7_16),
		.out_row (out_row_8_16),
		.out_col (out_col_8_16),
		.out_data (out_data_8_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_17;
	wire signed [DATA_WIDTH-1:0] out_col_8_17;
	wire signed [DATA_WIDTH-1:0] out_data_8_17;
	integer_mac_pe mac_pe_8_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_16),
		.in_col (out_col_7_17),
		.out_row (out_row_8_17),
		.out_col (out_col_8_17),
		.out_data (out_data_8_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_18;
	wire signed [DATA_WIDTH-1:0] out_col_8_18;
	wire signed [DATA_WIDTH-1:0] out_data_8_18;
	integer_mac_pe mac_pe_8_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_17),
		.in_col (out_col_7_18),
		.out_row (out_row_8_18),
		.out_col (out_col_8_18),
		.out_data (out_data_8_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_19;
	wire signed [DATA_WIDTH-1:0] out_col_8_19;
	wire signed [DATA_WIDTH-1:0] out_data_8_19;
	integer_mac_pe mac_pe_8_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_18),
		.in_col (out_col_7_19),
		.out_row (out_row_8_19),
		.out_col (out_col_8_19),
		.out_data (out_data_8_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_20;
	wire signed [DATA_WIDTH-1:0] out_col_8_20;
	wire signed [DATA_WIDTH-1:0] out_data_8_20;
	integer_mac_pe mac_pe_8_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_19),
		.in_col (out_col_7_20),
		.out_row (out_row_8_20),
		.out_col (out_col_8_20),
		.out_data (out_data_8_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_21;
	wire signed [DATA_WIDTH-1:0] out_col_8_21;
	wire signed [DATA_WIDTH-1:0] out_data_8_21;
	integer_mac_pe mac_pe_8_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_20),
		.in_col (out_col_7_21),
		.out_row (out_row_8_21),
		.out_col (out_col_8_21),
		.out_data (out_data_8_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_22;
	wire signed [DATA_WIDTH-1:0] out_col_8_22;
	wire signed [DATA_WIDTH-1:0] out_data_8_22;
	integer_mac_pe mac_pe_8_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_21),
		.in_col (out_col_7_22),
		.out_row (out_row_8_22),
		.out_col (out_col_8_22),
		.out_data (out_data_8_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_23;
	wire signed [DATA_WIDTH-1:0] out_col_8_23;
	wire signed [DATA_WIDTH-1:0] out_data_8_23;
	integer_mac_pe mac_pe_8_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_22),
		.in_col (out_col_7_23),
		.out_row (out_row_8_23),
		.out_col (out_col_8_23),
		.out_data (out_data_8_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_24;
	wire signed [DATA_WIDTH-1:0] out_col_8_24;
	wire signed [DATA_WIDTH-1:0] out_data_8_24;
	integer_mac_pe mac_pe_8_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_23),
		.in_col (out_col_7_24),
		.out_row (out_row_8_24),
		.out_col (out_col_8_24),
		.out_data (out_data_8_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_25;
	wire signed [DATA_WIDTH-1:0] out_col_8_25;
	wire signed [DATA_WIDTH-1:0] out_data_8_25;
	integer_mac_pe mac_pe_8_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_24),
		.in_col (out_col_7_25),
		.out_row (out_row_8_25),
		.out_col (out_col_8_25),
		.out_data (out_data_8_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_26;
	wire signed [DATA_WIDTH-1:0] out_col_8_26;
	wire signed [DATA_WIDTH-1:0] out_data_8_26;
	integer_mac_pe mac_pe_8_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_25),
		.in_col (out_col_7_26),
		.out_row (out_row_8_26),
		.out_col (out_col_8_26),
		.out_data (out_data_8_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_27;
	wire signed [DATA_WIDTH-1:0] out_col_8_27;
	wire signed [DATA_WIDTH-1:0] out_data_8_27;
	integer_mac_pe mac_pe_8_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_26),
		.in_col (out_col_7_27),
		.out_row (out_row_8_27),
		.out_col (out_col_8_27),
		.out_data (out_data_8_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_28;
	wire signed [DATA_WIDTH-1:0] out_col_8_28;
	wire signed [DATA_WIDTH-1:0] out_data_8_28;
	integer_mac_pe mac_pe_8_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_27),
		.in_col (out_col_7_28),
		.out_row (out_row_8_28),
		.out_col (out_col_8_28),
		.out_data (out_data_8_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_29;
	wire signed [DATA_WIDTH-1:0] out_col_8_29;
	wire signed [DATA_WIDTH-1:0] out_data_8_29;
	integer_mac_pe mac_pe_8_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_28),
		.in_col (out_col_7_29),
		.out_row (out_row_8_29),
		.out_col (out_col_8_29),
		.out_data (out_data_8_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_30;
	wire signed [DATA_WIDTH-1:0] out_col_8_30;
	wire signed [DATA_WIDTH-1:0] out_data_8_30;
	integer_mac_pe mac_pe_8_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_29),
		.in_col (out_col_7_30),
		.out_row (out_row_8_30),
		.out_col (out_col_8_30),
		.out_data (out_data_8_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_8_31;
	wire signed [DATA_WIDTH-1:0] out_col_8_31;
	wire signed [DATA_WIDTH-1:0] out_data_8_31;
	integer_mac_pe mac_pe_8_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_8_30),
		.in_col (out_col_7_31),
		.out_row (out_row_8_31),
		.out_col (out_col_8_31),
		.out_data (out_data_8_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_0;
	wire signed [DATA_WIDTH-1:0] out_col_9_0;
	wire signed [DATA_WIDTH-1:0] out_data_9_0;
	integer_mac_pe mac_pe_9_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_9_out),
		.in_col (out_col_8_0),
		.out_row (out_row_9_0),
		.out_col (out_col_9_0),
		.out_data (out_data_9_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_1;
	wire signed [DATA_WIDTH-1:0] out_col_9_1;
	wire signed [DATA_WIDTH-1:0] out_data_9_1;
	integer_mac_pe mac_pe_9_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_0),
		.in_col (out_col_8_1),
		.out_row (out_row_9_1),
		.out_col (out_col_9_1),
		.out_data (out_data_9_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_2;
	wire signed [DATA_WIDTH-1:0] out_col_9_2;
	wire signed [DATA_WIDTH-1:0] out_data_9_2;
	integer_mac_pe mac_pe_9_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_1),
		.in_col (out_col_8_2),
		.out_row (out_row_9_2),
		.out_col (out_col_9_2),
		.out_data (out_data_9_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_3;
	wire signed [DATA_WIDTH-1:0] out_col_9_3;
	wire signed [DATA_WIDTH-1:0] out_data_9_3;
	integer_mac_pe mac_pe_9_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_2),
		.in_col (out_col_8_3),
		.out_row (out_row_9_3),
		.out_col (out_col_9_3),
		.out_data (out_data_9_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_4;
	wire signed [DATA_WIDTH-1:0] out_col_9_4;
	wire signed [DATA_WIDTH-1:0] out_data_9_4;
	integer_mac_pe mac_pe_9_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_3),
		.in_col (out_col_8_4),
		.out_row (out_row_9_4),
		.out_col (out_col_9_4),
		.out_data (out_data_9_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_5;
	wire signed [DATA_WIDTH-1:0] out_col_9_5;
	wire signed [DATA_WIDTH-1:0] out_data_9_5;
	integer_mac_pe mac_pe_9_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_4),
		.in_col (out_col_8_5),
		.out_row (out_row_9_5),
		.out_col (out_col_9_5),
		.out_data (out_data_9_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_6;
	wire signed [DATA_WIDTH-1:0] out_col_9_6;
	wire signed [DATA_WIDTH-1:0] out_data_9_6;
	integer_mac_pe mac_pe_9_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_5),
		.in_col (out_col_8_6),
		.out_row (out_row_9_6),
		.out_col (out_col_9_6),
		.out_data (out_data_9_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_7;
	wire signed [DATA_WIDTH-1:0] out_col_9_7;
	wire signed [DATA_WIDTH-1:0] out_data_9_7;
	integer_mac_pe mac_pe_9_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_6),
		.in_col (out_col_8_7),
		.out_row (out_row_9_7),
		.out_col (out_col_9_7),
		.out_data (out_data_9_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_8;
	wire signed [DATA_WIDTH-1:0] out_col_9_8;
	wire signed [DATA_WIDTH-1:0] out_data_9_8;
	integer_mac_pe mac_pe_9_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_7),
		.in_col (out_col_8_8),
		.out_row (out_row_9_8),
		.out_col (out_col_9_8),
		.out_data (out_data_9_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_9;
	wire signed [DATA_WIDTH-1:0] out_col_9_9;
	wire signed [DATA_WIDTH-1:0] out_data_9_9;
	integer_mac_pe mac_pe_9_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_8),
		.in_col (out_col_8_9),
		.out_row (out_row_9_9),
		.out_col (out_col_9_9),
		.out_data (out_data_9_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_10;
	wire signed [DATA_WIDTH-1:0] out_col_9_10;
	wire signed [DATA_WIDTH-1:0] out_data_9_10;
	integer_mac_pe mac_pe_9_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_9),
		.in_col (out_col_8_10),
		.out_row (out_row_9_10),
		.out_col (out_col_9_10),
		.out_data (out_data_9_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_11;
	wire signed [DATA_WIDTH-1:0] out_col_9_11;
	wire signed [DATA_WIDTH-1:0] out_data_9_11;
	integer_mac_pe mac_pe_9_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_10),
		.in_col (out_col_8_11),
		.out_row (out_row_9_11),
		.out_col (out_col_9_11),
		.out_data (out_data_9_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_12;
	wire signed [DATA_WIDTH-1:0] out_col_9_12;
	wire signed [DATA_WIDTH-1:0] out_data_9_12;
	integer_mac_pe mac_pe_9_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_11),
		.in_col (out_col_8_12),
		.out_row (out_row_9_12),
		.out_col (out_col_9_12),
		.out_data (out_data_9_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_13;
	wire signed [DATA_WIDTH-1:0] out_col_9_13;
	wire signed [DATA_WIDTH-1:0] out_data_9_13;
	integer_mac_pe mac_pe_9_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_12),
		.in_col (out_col_8_13),
		.out_row (out_row_9_13),
		.out_col (out_col_9_13),
		.out_data (out_data_9_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_14;
	wire signed [DATA_WIDTH-1:0] out_col_9_14;
	wire signed [DATA_WIDTH-1:0] out_data_9_14;
	integer_mac_pe mac_pe_9_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_13),
		.in_col (out_col_8_14),
		.out_row (out_row_9_14),
		.out_col (out_col_9_14),
		.out_data (out_data_9_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_15;
	wire signed [DATA_WIDTH-1:0] out_col_9_15;
	wire signed [DATA_WIDTH-1:0] out_data_9_15;
	integer_mac_pe mac_pe_9_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_14),
		.in_col (out_col_8_15),
		.out_row (out_row_9_15),
		.out_col (out_col_9_15),
		.out_data (out_data_9_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_16;
	wire signed [DATA_WIDTH-1:0] out_col_9_16;
	wire signed [DATA_WIDTH-1:0] out_data_9_16;
	integer_mac_pe mac_pe_9_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_15),
		.in_col (out_col_8_16),
		.out_row (out_row_9_16),
		.out_col (out_col_9_16),
		.out_data (out_data_9_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_17;
	wire signed [DATA_WIDTH-1:0] out_col_9_17;
	wire signed [DATA_WIDTH-1:0] out_data_9_17;
	integer_mac_pe mac_pe_9_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_16),
		.in_col (out_col_8_17),
		.out_row (out_row_9_17),
		.out_col (out_col_9_17),
		.out_data (out_data_9_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_18;
	wire signed [DATA_WIDTH-1:0] out_col_9_18;
	wire signed [DATA_WIDTH-1:0] out_data_9_18;
	integer_mac_pe mac_pe_9_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_17),
		.in_col (out_col_8_18),
		.out_row (out_row_9_18),
		.out_col (out_col_9_18),
		.out_data (out_data_9_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_19;
	wire signed [DATA_WIDTH-1:0] out_col_9_19;
	wire signed [DATA_WIDTH-1:0] out_data_9_19;
	integer_mac_pe mac_pe_9_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_18),
		.in_col (out_col_8_19),
		.out_row (out_row_9_19),
		.out_col (out_col_9_19),
		.out_data (out_data_9_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_20;
	wire signed [DATA_WIDTH-1:0] out_col_9_20;
	wire signed [DATA_WIDTH-1:0] out_data_9_20;
	integer_mac_pe mac_pe_9_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_19),
		.in_col (out_col_8_20),
		.out_row (out_row_9_20),
		.out_col (out_col_9_20),
		.out_data (out_data_9_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_21;
	wire signed [DATA_WIDTH-1:0] out_col_9_21;
	wire signed [DATA_WIDTH-1:0] out_data_9_21;
	integer_mac_pe mac_pe_9_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_20),
		.in_col (out_col_8_21),
		.out_row (out_row_9_21),
		.out_col (out_col_9_21),
		.out_data (out_data_9_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_22;
	wire signed [DATA_WIDTH-1:0] out_col_9_22;
	wire signed [DATA_WIDTH-1:0] out_data_9_22;
	integer_mac_pe mac_pe_9_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_21),
		.in_col (out_col_8_22),
		.out_row (out_row_9_22),
		.out_col (out_col_9_22),
		.out_data (out_data_9_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_23;
	wire signed [DATA_WIDTH-1:0] out_col_9_23;
	wire signed [DATA_WIDTH-1:0] out_data_9_23;
	integer_mac_pe mac_pe_9_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_22),
		.in_col (out_col_8_23),
		.out_row (out_row_9_23),
		.out_col (out_col_9_23),
		.out_data (out_data_9_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_24;
	wire signed [DATA_WIDTH-1:0] out_col_9_24;
	wire signed [DATA_WIDTH-1:0] out_data_9_24;
	integer_mac_pe mac_pe_9_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_23),
		.in_col (out_col_8_24),
		.out_row (out_row_9_24),
		.out_col (out_col_9_24),
		.out_data (out_data_9_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_25;
	wire signed [DATA_WIDTH-1:0] out_col_9_25;
	wire signed [DATA_WIDTH-1:0] out_data_9_25;
	integer_mac_pe mac_pe_9_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_24),
		.in_col (out_col_8_25),
		.out_row (out_row_9_25),
		.out_col (out_col_9_25),
		.out_data (out_data_9_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_26;
	wire signed [DATA_WIDTH-1:0] out_col_9_26;
	wire signed [DATA_WIDTH-1:0] out_data_9_26;
	integer_mac_pe mac_pe_9_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_25),
		.in_col (out_col_8_26),
		.out_row (out_row_9_26),
		.out_col (out_col_9_26),
		.out_data (out_data_9_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_27;
	wire signed [DATA_WIDTH-1:0] out_col_9_27;
	wire signed [DATA_WIDTH-1:0] out_data_9_27;
	integer_mac_pe mac_pe_9_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_26),
		.in_col (out_col_8_27),
		.out_row (out_row_9_27),
		.out_col (out_col_9_27),
		.out_data (out_data_9_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_28;
	wire signed [DATA_WIDTH-1:0] out_col_9_28;
	wire signed [DATA_WIDTH-1:0] out_data_9_28;
	integer_mac_pe mac_pe_9_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_27),
		.in_col (out_col_8_28),
		.out_row (out_row_9_28),
		.out_col (out_col_9_28),
		.out_data (out_data_9_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_29;
	wire signed [DATA_WIDTH-1:0] out_col_9_29;
	wire signed [DATA_WIDTH-1:0] out_data_9_29;
	integer_mac_pe mac_pe_9_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_28),
		.in_col (out_col_8_29),
		.out_row (out_row_9_29),
		.out_col (out_col_9_29),
		.out_data (out_data_9_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_30;
	wire signed [DATA_WIDTH-1:0] out_col_9_30;
	wire signed [DATA_WIDTH-1:0] out_data_9_30;
	integer_mac_pe mac_pe_9_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_29),
		.in_col (out_col_8_30),
		.out_row (out_row_9_30),
		.out_col (out_col_9_30),
		.out_data (out_data_9_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_9_31;
	wire signed [DATA_WIDTH-1:0] out_col_9_31;
	wire signed [DATA_WIDTH-1:0] out_data_9_31;
	integer_mac_pe mac_pe_9_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_9_30),
		.in_col (out_col_8_31),
		.out_row (out_row_9_31),
		.out_col (out_col_9_31),
		.out_data (out_data_9_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_0;
	wire signed [DATA_WIDTH-1:0] out_col_10_0;
	wire signed [DATA_WIDTH-1:0] out_data_10_0;
	integer_mac_pe mac_pe_10_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_10_out),
		.in_col (out_col_9_0),
		.out_row (out_row_10_0),
		.out_col (out_col_10_0),
		.out_data (out_data_10_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_1;
	wire signed [DATA_WIDTH-1:0] out_col_10_1;
	wire signed [DATA_WIDTH-1:0] out_data_10_1;
	integer_mac_pe mac_pe_10_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_0),
		.in_col (out_col_9_1),
		.out_row (out_row_10_1),
		.out_col (out_col_10_1),
		.out_data (out_data_10_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_2;
	wire signed [DATA_WIDTH-1:0] out_col_10_2;
	wire signed [DATA_WIDTH-1:0] out_data_10_2;
	integer_mac_pe mac_pe_10_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_1),
		.in_col (out_col_9_2),
		.out_row (out_row_10_2),
		.out_col (out_col_10_2),
		.out_data (out_data_10_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_3;
	wire signed [DATA_WIDTH-1:0] out_col_10_3;
	wire signed [DATA_WIDTH-1:0] out_data_10_3;
	integer_mac_pe mac_pe_10_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_2),
		.in_col (out_col_9_3),
		.out_row (out_row_10_3),
		.out_col (out_col_10_3),
		.out_data (out_data_10_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_4;
	wire signed [DATA_WIDTH-1:0] out_col_10_4;
	wire signed [DATA_WIDTH-1:0] out_data_10_4;
	integer_mac_pe mac_pe_10_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_3),
		.in_col (out_col_9_4),
		.out_row (out_row_10_4),
		.out_col (out_col_10_4),
		.out_data (out_data_10_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_5;
	wire signed [DATA_WIDTH-1:0] out_col_10_5;
	wire signed [DATA_WIDTH-1:0] out_data_10_5;
	integer_mac_pe mac_pe_10_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_4),
		.in_col (out_col_9_5),
		.out_row (out_row_10_5),
		.out_col (out_col_10_5),
		.out_data (out_data_10_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_6;
	wire signed [DATA_WIDTH-1:0] out_col_10_6;
	wire signed [DATA_WIDTH-1:0] out_data_10_6;
	integer_mac_pe mac_pe_10_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_5),
		.in_col (out_col_9_6),
		.out_row (out_row_10_6),
		.out_col (out_col_10_6),
		.out_data (out_data_10_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_7;
	wire signed [DATA_WIDTH-1:0] out_col_10_7;
	wire signed [DATA_WIDTH-1:0] out_data_10_7;
	integer_mac_pe mac_pe_10_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_6),
		.in_col (out_col_9_7),
		.out_row (out_row_10_7),
		.out_col (out_col_10_7),
		.out_data (out_data_10_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_8;
	wire signed [DATA_WIDTH-1:0] out_col_10_8;
	wire signed [DATA_WIDTH-1:0] out_data_10_8;
	integer_mac_pe mac_pe_10_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_7),
		.in_col (out_col_9_8),
		.out_row (out_row_10_8),
		.out_col (out_col_10_8),
		.out_data (out_data_10_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_9;
	wire signed [DATA_WIDTH-1:0] out_col_10_9;
	wire signed [DATA_WIDTH-1:0] out_data_10_9;
	integer_mac_pe mac_pe_10_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_8),
		.in_col (out_col_9_9),
		.out_row (out_row_10_9),
		.out_col (out_col_10_9),
		.out_data (out_data_10_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_10;
	wire signed [DATA_WIDTH-1:0] out_col_10_10;
	wire signed [DATA_WIDTH-1:0] out_data_10_10;
	integer_mac_pe mac_pe_10_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_9),
		.in_col (out_col_9_10),
		.out_row (out_row_10_10),
		.out_col (out_col_10_10),
		.out_data (out_data_10_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_11;
	wire signed [DATA_WIDTH-1:0] out_col_10_11;
	wire signed [DATA_WIDTH-1:0] out_data_10_11;
	integer_mac_pe mac_pe_10_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_10),
		.in_col (out_col_9_11),
		.out_row (out_row_10_11),
		.out_col (out_col_10_11),
		.out_data (out_data_10_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_12;
	wire signed [DATA_WIDTH-1:0] out_col_10_12;
	wire signed [DATA_WIDTH-1:0] out_data_10_12;
	integer_mac_pe mac_pe_10_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_11),
		.in_col (out_col_9_12),
		.out_row (out_row_10_12),
		.out_col (out_col_10_12),
		.out_data (out_data_10_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_13;
	wire signed [DATA_WIDTH-1:0] out_col_10_13;
	wire signed [DATA_WIDTH-1:0] out_data_10_13;
	integer_mac_pe mac_pe_10_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_12),
		.in_col (out_col_9_13),
		.out_row (out_row_10_13),
		.out_col (out_col_10_13),
		.out_data (out_data_10_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_14;
	wire signed [DATA_WIDTH-1:0] out_col_10_14;
	wire signed [DATA_WIDTH-1:0] out_data_10_14;
	integer_mac_pe mac_pe_10_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_13),
		.in_col (out_col_9_14),
		.out_row (out_row_10_14),
		.out_col (out_col_10_14),
		.out_data (out_data_10_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_15;
	wire signed [DATA_WIDTH-1:0] out_col_10_15;
	wire signed [DATA_WIDTH-1:0] out_data_10_15;
	integer_mac_pe mac_pe_10_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_14),
		.in_col (out_col_9_15),
		.out_row (out_row_10_15),
		.out_col (out_col_10_15),
		.out_data (out_data_10_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_16;
	wire signed [DATA_WIDTH-1:0] out_col_10_16;
	wire signed [DATA_WIDTH-1:0] out_data_10_16;
	integer_mac_pe mac_pe_10_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_15),
		.in_col (out_col_9_16),
		.out_row (out_row_10_16),
		.out_col (out_col_10_16),
		.out_data (out_data_10_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_17;
	wire signed [DATA_WIDTH-1:0] out_col_10_17;
	wire signed [DATA_WIDTH-1:0] out_data_10_17;
	integer_mac_pe mac_pe_10_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_16),
		.in_col (out_col_9_17),
		.out_row (out_row_10_17),
		.out_col (out_col_10_17),
		.out_data (out_data_10_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_18;
	wire signed [DATA_WIDTH-1:0] out_col_10_18;
	wire signed [DATA_WIDTH-1:0] out_data_10_18;
	integer_mac_pe mac_pe_10_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_17),
		.in_col (out_col_9_18),
		.out_row (out_row_10_18),
		.out_col (out_col_10_18),
		.out_data (out_data_10_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_19;
	wire signed [DATA_WIDTH-1:0] out_col_10_19;
	wire signed [DATA_WIDTH-1:0] out_data_10_19;
	integer_mac_pe mac_pe_10_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_18),
		.in_col (out_col_9_19),
		.out_row (out_row_10_19),
		.out_col (out_col_10_19),
		.out_data (out_data_10_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_20;
	wire signed [DATA_WIDTH-1:0] out_col_10_20;
	wire signed [DATA_WIDTH-1:0] out_data_10_20;
	integer_mac_pe mac_pe_10_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_19),
		.in_col (out_col_9_20),
		.out_row (out_row_10_20),
		.out_col (out_col_10_20),
		.out_data (out_data_10_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_21;
	wire signed [DATA_WIDTH-1:0] out_col_10_21;
	wire signed [DATA_WIDTH-1:0] out_data_10_21;
	integer_mac_pe mac_pe_10_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_20),
		.in_col (out_col_9_21),
		.out_row (out_row_10_21),
		.out_col (out_col_10_21),
		.out_data (out_data_10_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_22;
	wire signed [DATA_WIDTH-1:0] out_col_10_22;
	wire signed [DATA_WIDTH-1:0] out_data_10_22;
	integer_mac_pe mac_pe_10_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_21),
		.in_col (out_col_9_22),
		.out_row (out_row_10_22),
		.out_col (out_col_10_22),
		.out_data (out_data_10_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_23;
	wire signed [DATA_WIDTH-1:0] out_col_10_23;
	wire signed [DATA_WIDTH-1:0] out_data_10_23;
	integer_mac_pe mac_pe_10_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_22),
		.in_col (out_col_9_23),
		.out_row (out_row_10_23),
		.out_col (out_col_10_23),
		.out_data (out_data_10_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_24;
	wire signed [DATA_WIDTH-1:0] out_col_10_24;
	wire signed [DATA_WIDTH-1:0] out_data_10_24;
	integer_mac_pe mac_pe_10_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_23),
		.in_col (out_col_9_24),
		.out_row (out_row_10_24),
		.out_col (out_col_10_24),
		.out_data (out_data_10_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_25;
	wire signed [DATA_WIDTH-1:0] out_col_10_25;
	wire signed [DATA_WIDTH-1:0] out_data_10_25;
	integer_mac_pe mac_pe_10_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_24),
		.in_col (out_col_9_25),
		.out_row (out_row_10_25),
		.out_col (out_col_10_25),
		.out_data (out_data_10_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_26;
	wire signed [DATA_WIDTH-1:0] out_col_10_26;
	wire signed [DATA_WIDTH-1:0] out_data_10_26;
	integer_mac_pe mac_pe_10_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_25),
		.in_col (out_col_9_26),
		.out_row (out_row_10_26),
		.out_col (out_col_10_26),
		.out_data (out_data_10_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_27;
	wire signed [DATA_WIDTH-1:0] out_col_10_27;
	wire signed [DATA_WIDTH-1:0] out_data_10_27;
	integer_mac_pe mac_pe_10_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_26),
		.in_col (out_col_9_27),
		.out_row (out_row_10_27),
		.out_col (out_col_10_27),
		.out_data (out_data_10_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_28;
	wire signed [DATA_WIDTH-1:0] out_col_10_28;
	wire signed [DATA_WIDTH-1:0] out_data_10_28;
	integer_mac_pe mac_pe_10_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_27),
		.in_col (out_col_9_28),
		.out_row (out_row_10_28),
		.out_col (out_col_10_28),
		.out_data (out_data_10_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_29;
	wire signed [DATA_WIDTH-1:0] out_col_10_29;
	wire signed [DATA_WIDTH-1:0] out_data_10_29;
	integer_mac_pe mac_pe_10_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_28),
		.in_col (out_col_9_29),
		.out_row (out_row_10_29),
		.out_col (out_col_10_29),
		.out_data (out_data_10_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_30;
	wire signed [DATA_WIDTH-1:0] out_col_10_30;
	wire signed [DATA_WIDTH-1:0] out_data_10_30;
	integer_mac_pe mac_pe_10_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_29),
		.in_col (out_col_9_30),
		.out_row (out_row_10_30),
		.out_col (out_col_10_30),
		.out_data (out_data_10_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_10_31;
	wire signed [DATA_WIDTH-1:0] out_col_10_31;
	wire signed [DATA_WIDTH-1:0] out_data_10_31;
	integer_mac_pe mac_pe_10_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_10_30),
		.in_col (out_col_9_31),
		.out_row (out_row_10_31),
		.out_col (out_col_10_31),
		.out_data (out_data_10_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_0;
	wire signed [DATA_WIDTH-1:0] out_col_11_0;
	wire signed [DATA_WIDTH-1:0] out_data_11_0;
	integer_mac_pe mac_pe_11_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_11_out),
		.in_col (out_col_10_0),
		.out_row (out_row_11_0),
		.out_col (out_col_11_0),
		.out_data (out_data_11_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_1;
	wire signed [DATA_WIDTH-1:0] out_col_11_1;
	wire signed [DATA_WIDTH-1:0] out_data_11_1;
	integer_mac_pe mac_pe_11_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_0),
		.in_col (out_col_10_1),
		.out_row (out_row_11_1),
		.out_col (out_col_11_1),
		.out_data (out_data_11_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_2;
	wire signed [DATA_WIDTH-1:0] out_col_11_2;
	wire signed [DATA_WIDTH-1:0] out_data_11_2;
	integer_mac_pe mac_pe_11_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_1),
		.in_col (out_col_10_2),
		.out_row (out_row_11_2),
		.out_col (out_col_11_2),
		.out_data (out_data_11_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_3;
	wire signed [DATA_WIDTH-1:0] out_col_11_3;
	wire signed [DATA_WIDTH-1:0] out_data_11_3;
	integer_mac_pe mac_pe_11_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_2),
		.in_col (out_col_10_3),
		.out_row (out_row_11_3),
		.out_col (out_col_11_3),
		.out_data (out_data_11_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_4;
	wire signed [DATA_WIDTH-1:0] out_col_11_4;
	wire signed [DATA_WIDTH-1:0] out_data_11_4;
	integer_mac_pe mac_pe_11_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_3),
		.in_col (out_col_10_4),
		.out_row (out_row_11_4),
		.out_col (out_col_11_4),
		.out_data (out_data_11_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_5;
	wire signed [DATA_WIDTH-1:0] out_col_11_5;
	wire signed [DATA_WIDTH-1:0] out_data_11_5;
	integer_mac_pe mac_pe_11_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_4),
		.in_col (out_col_10_5),
		.out_row (out_row_11_5),
		.out_col (out_col_11_5),
		.out_data (out_data_11_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_6;
	wire signed [DATA_WIDTH-1:0] out_col_11_6;
	wire signed [DATA_WIDTH-1:0] out_data_11_6;
	integer_mac_pe mac_pe_11_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_5),
		.in_col (out_col_10_6),
		.out_row (out_row_11_6),
		.out_col (out_col_11_6),
		.out_data (out_data_11_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_7;
	wire signed [DATA_WIDTH-1:0] out_col_11_7;
	wire signed [DATA_WIDTH-1:0] out_data_11_7;
	integer_mac_pe mac_pe_11_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_6),
		.in_col (out_col_10_7),
		.out_row (out_row_11_7),
		.out_col (out_col_11_7),
		.out_data (out_data_11_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_8;
	wire signed [DATA_WIDTH-1:0] out_col_11_8;
	wire signed [DATA_WIDTH-1:0] out_data_11_8;
	integer_mac_pe mac_pe_11_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_7),
		.in_col (out_col_10_8),
		.out_row (out_row_11_8),
		.out_col (out_col_11_8),
		.out_data (out_data_11_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_9;
	wire signed [DATA_WIDTH-1:0] out_col_11_9;
	wire signed [DATA_WIDTH-1:0] out_data_11_9;
	integer_mac_pe mac_pe_11_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_8),
		.in_col (out_col_10_9),
		.out_row (out_row_11_9),
		.out_col (out_col_11_9),
		.out_data (out_data_11_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_10;
	wire signed [DATA_WIDTH-1:0] out_col_11_10;
	wire signed [DATA_WIDTH-1:0] out_data_11_10;
	integer_mac_pe mac_pe_11_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_9),
		.in_col (out_col_10_10),
		.out_row (out_row_11_10),
		.out_col (out_col_11_10),
		.out_data (out_data_11_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_11;
	wire signed [DATA_WIDTH-1:0] out_col_11_11;
	wire signed [DATA_WIDTH-1:0] out_data_11_11;
	integer_mac_pe mac_pe_11_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_10),
		.in_col (out_col_10_11),
		.out_row (out_row_11_11),
		.out_col (out_col_11_11),
		.out_data (out_data_11_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_12;
	wire signed [DATA_WIDTH-1:0] out_col_11_12;
	wire signed [DATA_WIDTH-1:0] out_data_11_12;
	integer_mac_pe mac_pe_11_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_11),
		.in_col (out_col_10_12),
		.out_row (out_row_11_12),
		.out_col (out_col_11_12),
		.out_data (out_data_11_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_13;
	wire signed [DATA_WIDTH-1:0] out_col_11_13;
	wire signed [DATA_WIDTH-1:0] out_data_11_13;
	integer_mac_pe mac_pe_11_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_12),
		.in_col (out_col_10_13),
		.out_row (out_row_11_13),
		.out_col (out_col_11_13),
		.out_data (out_data_11_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_14;
	wire signed [DATA_WIDTH-1:0] out_col_11_14;
	wire signed [DATA_WIDTH-1:0] out_data_11_14;
	integer_mac_pe mac_pe_11_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_13),
		.in_col (out_col_10_14),
		.out_row (out_row_11_14),
		.out_col (out_col_11_14),
		.out_data (out_data_11_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_15;
	wire signed [DATA_WIDTH-1:0] out_col_11_15;
	wire signed [DATA_WIDTH-1:0] out_data_11_15;
	integer_mac_pe mac_pe_11_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_14),
		.in_col (out_col_10_15),
		.out_row (out_row_11_15),
		.out_col (out_col_11_15),
		.out_data (out_data_11_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_16;
	wire signed [DATA_WIDTH-1:0] out_col_11_16;
	wire signed [DATA_WIDTH-1:0] out_data_11_16;
	integer_mac_pe mac_pe_11_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_15),
		.in_col (out_col_10_16),
		.out_row (out_row_11_16),
		.out_col (out_col_11_16),
		.out_data (out_data_11_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_17;
	wire signed [DATA_WIDTH-1:0] out_col_11_17;
	wire signed [DATA_WIDTH-1:0] out_data_11_17;
	integer_mac_pe mac_pe_11_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_16),
		.in_col (out_col_10_17),
		.out_row (out_row_11_17),
		.out_col (out_col_11_17),
		.out_data (out_data_11_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_18;
	wire signed [DATA_WIDTH-1:0] out_col_11_18;
	wire signed [DATA_WIDTH-1:0] out_data_11_18;
	integer_mac_pe mac_pe_11_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_17),
		.in_col (out_col_10_18),
		.out_row (out_row_11_18),
		.out_col (out_col_11_18),
		.out_data (out_data_11_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_19;
	wire signed [DATA_WIDTH-1:0] out_col_11_19;
	wire signed [DATA_WIDTH-1:0] out_data_11_19;
	integer_mac_pe mac_pe_11_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_18),
		.in_col (out_col_10_19),
		.out_row (out_row_11_19),
		.out_col (out_col_11_19),
		.out_data (out_data_11_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_20;
	wire signed [DATA_WIDTH-1:0] out_col_11_20;
	wire signed [DATA_WIDTH-1:0] out_data_11_20;
	integer_mac_pe mac_pe_11_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_19),
		.in_col (out_col_10_20),
		.out_row (out_row_11_20),
		.out_col (out_col_11_20),
		.out_data (out_data_11_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_21;
	wire signed [DATA_WIDTH-1:0] out_col_11_21;
	wire signed [DATA_WIDTH-1:0] out_data_11_21;
	integer_mac_pe mac_pe_11_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_20),
		.in_col (out_col_10_21),
		.out_row (out_row_11_21),
		.out_col (out_col_11_21),
		.out_data (out_data_11_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_22;
	wire signed [DATA_WIDTH-1:0] out_col_11_22;
	wire signed [DATA_WIDTH-1:0] out_data_11_22;
	integer_mac_pe mac_pe_11_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_21),
		.in_col (out_col_10_22),
		.out_row (out_row_11_22),
		.out_col (out_col_11_22),
		.out_data (out_data_11_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_23;
	wire signed [DATA_WIDTH-1:0] out_col_11_23;
	wire signed [DATA_WIDTH-1:0] out_data_11_23;
	integer_mac_pe mac_pe_11_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_22),
		.in_col (out_col_10_23),
		.out_row (out_row_11_23),
		.out_col (out_col_11_23),
		.out_data (out_data_11_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_24;
	wire signed [DATA_WIDTH-1:0] out_col_11_24;
	wire signed [DATA_WIDTH-1:0] out_data_11_24;
	integer_mac_pe mac_pe_11_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_23),
		.in_col (out_col_10_24),
		.out_row (out_row_11_24),
		.out_col (out_col_11_24),
		.out_data (out_data_11_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_25;
	wire signed [DATA_WIDTH-1:0] out_col_11_25;
	wire signed [DATA_WIDTH-1:0] out_data_11_25;
	integer_mac_pe mac_pe_11_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_24),
		.in_col (out_col_10_25),
		.out_row (out_row_11_25),
		.out_col (out_col_11_25),
		.out_data (out_data_11_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_26;
	wire signed [DATA_WIDTH-1:0] out_col_11_26;
	wire signed [DATA_WIDTH-1:0] out_data_11_26;
	integer_mac_pe mac_pe_11_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_25),
		.in_col (out_col_10_26),
		.out_row (out_row_11_26),
		.out_col (out_col_11_26),
		.out_data (out_data_11_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_27;
	wire signed [DATA_WIDTH-1:0] out_col_11_27;
	wire signed [DATA_WIDTH-1:0] out_data_11_27;
	integer_mac_pe mac_pe_11_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_26),
		.in_col (out_col_10_27),
		.out_row (out_row_11_27),
		.out_col (out_col_11_27),
		.out_data (out_data_11_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_28;
	wire signed [DATA_WIDTH-1:0] out_col_11_28;
	wire signed [DATA_WIDTH-1:0] out_data_11_28;
	integer_mac_pe mac_pe_11_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_27),
		.in_col (out_col_10_28),
		.out_row (out_row_11_28),
		.out_col (out_col_11_28),
		.out_data (out_data_11_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_29;
	wire signed [DATA_WIDTH-1:0] out_col_11_29;
	wire signed [DATA_WIDTH-1:0] out_data_11_29;
	integer_mac_pe mac_pe_11_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_28),
		.in_col (out_col_10_29),
		.out_row (out_row_11_29),
		.out_col (out_col_11_29),
		.out_data (out_data_11_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_30;
	wire signed [DATA_WIDTH-1:0] out_col_11_30;
	wire signed [DATA_WIDTH-1:0] out_data_11_30;
	integer_mac_pe mac_pe_11_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_29),
		.in_col (out_col_10_30),
		.out_row (out_row_11_30),
		.out_col (out_col_11_30),
		.out_data (out_data_11_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_11_31;
	wire signed [DATA_WIDTH-1:0] out_col_11_31;
	wire signed [DATA_WIDTH-1:0] out_data_11_31;
	integer_mac_pe mac_pe_11_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_11_30),
		.in_col (out_col_10_31),
		.out_row (out_row_11_31),
		.out_col (out_col_11_31),
		.out_data (out_data_11_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_0;
	wire signed [DATA_WIDTH-1:0] out_col_12_0;
	wire signed [DATA_WIDTH-1:0] out_data_12_0;
	integer_mac_pe mac_pe_12_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_12_out),
		.in_col (out_col_11_0),
		.out_row (out_row_12_0),
		.out_col (out_col_12_0),
		.out_data (out_data_12_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_1;
	wire signed [DATA_WIDTH-1:0] out_col_12_1;
	wire signed [DATA_WIDTH-1:0] out_data_12_1;
	integer_mac_pe mac_pe_12_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_0),
		.in_col (out_col_11_1),
		.out_row (out_row_12_1),
		.out_col (out_col_12_1),
		.out_data (out_data_12_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_2;
	wire signed [DATA_WIDTH-1:0] out_col_12_2;
	wire signed [DATA_WIDTH-1:0] out_data_12_2;
	integer_mac_pe mac_pe_12_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_1),
		.in_col (out_col_11_2),
		.out_row (out_row_12_2),
		.out_col (out_col_12_2),
		.out_data (out_data_12_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_3;
	wire signed [DATA_WIDTH-1:0] out_col_12_3;
	wire signed [DATA_WIDTH-1:0] out_data_12_3;
	integer_mac_pe mac_pe_12_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_2),
		.in_col (out_col_11_3),
		.out_row (out_row_12_3),
		.out_col (out_col_12_3),
		.out_data (out_data_12_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_4;
	wire signed [DATA_WIDTH-1:0] out_col_12_4;
	wire signed [DATA_WIDTH-1:0] out_data_12_4;
	integer_mac_pe mac_pe_12_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_3),
		.in_col (out_col_11_4),
		.out_row (out_row_12_4),
		.out_col (out_col_12_4),
		.out_data (out_data_12_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_5;
	wire signed [DATA_WIDTH-1:0] out_col_12_5;
	wire signed [DATA_WIDTH-1:0] out_data_12_5;
	integer_mac_pe mac_pe_12_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_4),
		.in_col (out_col_11_5),
		.out_row (out_row_12_5),
		.out_col (out_col_12_5),
		.out_data (out_data_12_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_6;
	wire signed [DATA_WIDTH-1:0] out_col_12_6;
	wire signed [DATA_WIDTH-1:0] out_data_12_6;
	integer_mac_pe mac_pe_12_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_5),
		.in_col (out_col_11_6),
		.out_row (out_row_12_6),
		.out_col (out_col_12_6),
		.out_data (out_data_12_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_7;
	wire signed [DATA_WIDTH-1:0] out_col_12_7;
	wire signed [DATA_WIDTH-1:0] out_data_12_7;
	integer_mac_pe mac_pe_12_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_6),
		.in_col (out_col_11_7),
		.out_row (out_row_12_7),
		.out_col (out_col_12_7),
		.out_data (out_data_12_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_8;
	wire signed [DATA_WIDTH-1:0] out_col_12_8;
	wire signed [DATA_WIDTH-1:0] out_data_12_8;
	integer_mac_pe mac_pe_12_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_7),
		.in_col (out_col_11_8),
		.out_row (out_row_12_8),
		.out_col (out_col_12_8),
		.out_data (out_data_12_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_9;
	wire signed [DATA_WIDTH-1:0] out_col_12_9;
	wire signed [DATA_WIDTH-1:0] out_data_12_9;
	integer_mac_pe mac_pe_12_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_8),
		.in_col (out_col_11_9),
		.out_row (out_row_12_9),
		.out_col (out_col_12_9),
		.out_data (out_data_12_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_10;
	wire signed [DATA_WIDTH-1:0] out_col_12_10;
	wire signed [DATA_WIDTH-1:0] out_data_12_10;
	integer_mac_pe mac_pe_12_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_9),
		.in_col (out_col_11_10),
		.out_row (out_row_12_10),
		.out_col (out_col_12_10),
		.out_data (out_data_12_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_11;
	wire signed [DATA_WIDTH-1:0] out_col_12_11;
	wire signed [DATA_WIDTH-1:0] out_data_12_11;
	integer_mac_pe mac_pe_12_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_10),
		.in_col (out_col_11_11),
		.out_row (out_row_12_11),
		.out_col (out_col_12_11),
		.out_data (out_data_12_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_12;
	wire signed [DATA_WIDTH-1:0] out_col_12_12;
	wire signed [DATA_WIDTH-1:0] out_data_12_12;
	integer_mac_pe mac_pe_12_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_11),
		.in_col (out_col_11_12),
		.out_row (out_row_12_12),
		.out_col (out_col_12_12),
		.out_data (out_data_12_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_13;
	wire signed [DATA_WIDTH-1:0] out_col_12_13;
	wire signed [DATA_WIDTH-1:0] out_data_12_13;
	integer_mac_pe mac_pe_12_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_12),
		.in_col (out_col_11_13),
		.out_row (out_row_12_13),
		.out_col (out_col_12_13),
		.out_data (out_data_12_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_14;
	wire signed [DATA_WIDTH-1:0] out_col_12_14;
	wire signed [DATA_WIDTH-1:0] out_data_12_14;
	integer_mac_pe mac_pe_12_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_13),
		.in_col (out_col_11_14),
		.out_row (out_row_12_14),
		.out_col (out_col_12_14),
		.out_data (out_data_12_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_15;
	wire signed [DATA_WIDTH-1:0] out_col_12_15;
	wire signed [DATA_WIDTH-1:0] out_data_12_15;
	integer_mac_pe mac_pe_12_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_14),
		.in_col (out_col_11_15),
		.out_row (out_row_12_15),
		.out_col (out_col_12_15),
		.out_data (out_data_12_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_16;
	wire signed [DATA_WIDTH-1:0] out_col_12_16;
	wire signed [DATA_WIDTH-1:0] out_data_12_16;
	integer_mac_pe mac_pe_12_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_15),
		.in_col (out_col_11_16),
		.out_row (out_row_12_16),
		.out_col (out_col_12_16),
		.out_data (out_data_12_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_17;
	wire signed [DATA_WIDTH-1:0] out_col_12_17;
	wire signed [DATA_WIDTH-1:0] out_data_12_17;
	integer_mac_pe mac_pe_12_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_16),
		.in_col (out_col_11_17),
		.out_row (out_row_12_17),
		.out_col (out_col_12_17),
		.out_data (out_data_12_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_18;
	wire signed [DATA_WIDTH-1:0] out_col_12_18;
	wire signed [DATA_WIDTH-1:0] out_data_12_18;
	integer_mac_pe mac_pe_12_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_17),
		.in_col (out_col_11_18),
		.out_row (out_row_12_18),
		.out_col (out_col_12_18),
		.out_data (out_data_12_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_19;
	wire signed [DATA_WIDTH-1:0] out_col_12_19;
	wire signed [DATA_WIDTH-1:0] out_data_12_19;
	integer_mac_pe mac_pe_12_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_18),
		.in_col (out_col_11_19),
		.out_row (out_row_12_19),
		.out_col (out_col_12_19),
		.out_data (out_data_12_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_20;
	wire signed [DATA_WIDTH-1:0] out_col_12_20;
	wire signed [DATA_WIDTH-1:0] out_data_12_20;
	integer_mac_pe mac_pe_12_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_19),
		.in_col (out_col_11_20),
		.out_row (out_row_12_20),
		.out_col (out_col_12_20),
		.out_data (out_data_12_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_21;
	wire signed [DATA_WIDTH-1:0] out_col_12_21;
	wire signed [DATA_WIDTH-1:0] out_data_12_21;
	integer_mac_pe mac_pe_12_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_20),
		.in_col (out_col_11_21),
		.out_row (out_row_12_21),
		.out_col (out_col_12_21),
		.out_data (out_data_12_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_22;
	wire signed [DATA_WIDTH-1:0] out_col_12_22;
	wire signed [DATA_WIDTH-1:0] out_data_12_22;
	integer_mac_pe mac_pe_12_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_21),
		.in_col (out_col_11_22),
		.out_row (out_row_12_22),
		.out_col (out_col_12_22),
		.out_data (out_data_12_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_23;
	wire signed [DATA_WIDTH-1:0] out_col_12_23;
	wire signed [DATA_WIDTH-1:0] out_data_12_23;
	integer_mac_pe mac_pe_12_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_22),
		.in_col (out_col_11_23),
		.out_row (out_row_12_23),
		.out_col (out_col_12_23),
		.out_data (out_data_12_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_24;
	wire signed [DATA_WIDTH-1:0] out_col_12_24;
	wire signed [DATA_WIDTH-1:0] out_data_12_24;
	integer_mac_pe mac_pe_12_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_23),
		.in_col (out_col_11_24),
		.out_row (out_row_12_24),
		.out_col (out_col_12_24),
		.out_data (out_data_12_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_25;
	wire signed [DATA_WIDTH-1:0] out_col_12_25;
	wire signed [DATA_WIDTH-1:0] out_data_12_25;
	integer_mac_pe mac_pe_12_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_24),
		.in_col (out_col_11_25),
		.out_row (out_row_12_25),
		.out_col (out_col_12_25),
		.out_data (out_data_12_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_26;
	wire signed [DATA_WIDTH-1:0] out_col_12_26;
	wire signed [DATA_WIDTH-1:0] out_data_12_26;
	integer_mac_pe mac_pe_12_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_25),
		.in_col (out_col_11_26),
		.out_row (out_row_12_26),
		.out_col (out_col_12_26),
		.out_data (out_data_12_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_27;
	wire signed [DATA_WIDTH-1:0] out_col_12_27;
	wire signed [DATA_WIDTH-1:0] out_data_12_27;
	integer_mac_pe mac_pe_12_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_26),
		.in_col (out_col_11_27),
		.out_row (out_row_12_27),
		.out_col (out_col_12_27),
		.out_data (out_data_12_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_28;
	wire signed [DATA_WIDTH-1:0] out_col_12_28;
	wire signed [DATA_WIDTH-1:0] out_data_12_28;
	integer_mac_pe mac_pe_12_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_27),
		.in_col (out_col_11_28),
		.out_row (out_row_12_28),
		.out_col (out_col_12_28),
		.out_data (out_data_12_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_29;
	wire signed [DATA_WIDTH-1:0] out_col_12_29;
	wire signed [DATA_WIDTH-1:0] out_data_12_29;
	integer_mac_pe mac_pe_12_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_28),
		.in_col (out_col_11_29),
		.out_row (out_row_12_29),
		.out_col (out_col_12_29),
		.out_data (out_data_12_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_30;
	wire signed [DATA_WIDTH-1:0] out_col_12_30;
	wire signed [DATA_WIDTH-1:0] out_data_12_30;
	integer_mac_pe mac_pe_12_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_29),
		.in_col (out_col_11_30),
		.out_row (out_row_12_30),
		.out_col (out_col_12_30),
		.out_data (out_data_12_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_12_31;
	wire signed [DATA_WIDTH-1:0] out_col_12_31;
	wire signed [DATA_WIDTH-1:0] out_data_12_31;
	integer_mac_pe mac_pe_12_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_12_30),
		.in_col (out_col_11_31),
		.out_row (out_row_12_31),
		.out_col (out_col_12_31),
		.out_data (out_data_12_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_0;
	wire signed [DATA_WIDTH-1:0] out_col_13_0;
	wire signed [DATA_WIDTH-1:0] out_data_13_0;
	integer_mac_pe mac_pe_13_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_13_out),
		.in_col (out_col_12_0),
		.out_row (out_row_13_0),
		.out_col (out_col_13_0),
		.out_data (out_data_13_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_1;
	wire signed [DATA_WIDTH-1:0] out_col_13_1;
	wire signed [DATA_WIDTH-1:0] out_data_13_1;
	integer_mac_pe mac_pe_13_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_0),
		.in_col (out_col_12_1),
		.out_row (out_row_13_1),
		.out_col (out_col_13_1),
		.out_data (out_data_13_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_2;
	wire signed [DATA_WIDTH-1:0] out_col_13_2;
	wire signed [DATA_WIDTH-1:0] out_data_13_2;
	integer_mac_pe mac_pe_13_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_1),
		.in_col (out_col_12_2),
		.out_row (out_row_13_2),
		.out_col (out_col_13_2),
		.out_data (out_data_13_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_3;
	wire signed [DATA_WIDTH-1:0] out_col_13_3;
	wire signed [DATA_WIDTH-1:0] out_data_13_3;
	integer_mac_pe mac_pe_13_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_2),
		.in_col (out_col_12_3),
		.out_row (out_row_13_3),
		.out_col (out_col_13_3),
		.out_data (out_data_13_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_4;
	wire signed [DATA_WIDTH-1:0] out_col_13_4;
	wire signed [DATA_WIDTH-1:0] out_data_13_4;
	integer_mac_pe mac_pe_13_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_3),
		.in_col (out_col_12_4),
		.out_row (out_row_13_4),
		.out_col (out_col_13_4),
		.out_data (out_data_13_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_5;
	wire signed [DATA_WIDTH-1:0] out_col_13_5;
	wire signed [DATA_WIDTH-1:0] out_data_13_5;
	integer_mac_pe mac_pe_13_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_4),
		.in_col (out_col_12_5),
		.out_row (out_row_13_5),
		.out_col (out_col_13_5),
		.out_data (out_data_13_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_6;
	wire signed [DATA_WIDTH-1:0] out_col_13_6;
	wire signed [DATA_WIDTH-1:0] out_data_13_6;
	integer_mac_pe mac_pe_13_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_5),
		.in_col (out_col_12_6),
		.out_row (out_row_13_6),
		.out_col (out_col_13_6),
		.out_data (out_data_13_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_7;
	wire signed [DATA_WIDTH-1:0] out_col_13_7;
	wire signed [DATA_WIDTH-1:0] out_data_13_7;
	integer_mac_pe mac_pe_13_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_6),
		.in_col (out_col_12_7),
		.out_row (out_row_13_7),
		.out_col (out_col_13_7),
		.out_data (out_data_13_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_8;
	wire signed [DATA_WIDTH-1:0] out_col_13_8;
	wire signed [DATA_WIDTH-1:0] out_data_13_8;
	integer_mac_pe mac_pe_13_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_7),
		.in_col (out_col_12_8),
		.out_row (out_row_13_8),
		.out_col (out_col_13_8),
		.out_data (out_data_13_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_9;
	wire signed [DATA_WIDTH-1:0] out_col_13_9;
	wire signed [DATA_WIDTH-1:0] out_data_13_9;
	integer_mac_pe mac_pe_13_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_8),
		.in_col (out_col_12_9),
		.out_row (out_row_13_9),
		.out_col (out_col_13_9),
		.out_data (out_data_13_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_10;
	wire signed [DATA_WIDTH-1:0] out_col_13_10;
	wire signed [DATA_WIDTH-1:0] out_data_13_10;
	integer_mac_pe mac_pe_13_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_9),
		.in_col (out_col_12_10),
		.out_row (out_row_13_10),
		.out_col (out_col_13_10),
		.out_data (out_data_13_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_11;
	wire signed [DATA_WIDTH-1:0] out_col_13_11;
	wire signed [DATA_WIDTH-1:0] out_data_13_11;
	integer_mac_pe mac_pe_13_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_10),
		.in_col (out_col_12_11),
		.out_row (out_row_13_11),
		.out_col (out_col_13_11),
		.out_data (out_data_13_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_12;
	wire signed [DATA_WIDTH-1:0] out_col_13_12;
	wire signed [DATA_WIDTH-1:0] out_data_13_12;
	integer_mac_pe mac_pe_13_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_11),
		.in_col (out_col_12_12),
		.out_row (out_row_13_12),
		.out_col (out_col_13_12),
		.out_data (out_data_13_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_13;
	wire signed [DATA_WIDTH-1:0] out_col_13_13;
	wire signed [DATA_WIDTH-1:0] out_data_13_13;
	integer_mac_pe mac_pe_13_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_12),
		.in_col (out_col_12_13),
		.out_row (out_row_13_13),
		.out_col (out_col_13_13),
		.out_data (out_data_13_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_14;
	wire signed [DATA_WIDTH-1:0] out_col_13_14;
	wire signed [DATA_WIDTH-1:0] out_data_13_14;
	integer_mac_pe mac_pe_13_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_13),
		.in_col (out_col_12_14),
		.out_row (out_row_13_14),
		.out_col (out_col_13_14),
		.out_data (out_data_13_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_15;
	wire signed [DATA_WIDTH-1:0] out_col_13_15;
	wire signed [DATA_WIDTH-1:0] out_data_13_15;
	integer_mac_pe mac_pe_13_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_14),
		.in_col (out_col_12_15),
		.out_row (out_row_13_15),
		.out_col (out_col_13_15),
		.out_data (out_data_13_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_16;
	wire signed [DATA_WIDTH-1:0] out_col_13_16;
	wire signed [DATA_WIDTH-1:0] out_data_13_16;
	integer_mac_pe mac_pe_13_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_15),
		.in_col (out_col_12_16),
		.out_row (out_row_13_16),
		.out_col (out_col_13_16),
		.out_data (out_data_13_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_17;
	wire signed [DATA_WIDTH-1:0] out_col_13_17;
	wire signed [DATA_WIDTH-1:0] out_data_13_17;
	integer_mac_pe mac_pe_13_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_16),
		.in_col (out_col_12_17),
		.out_row (out_row_13_17),
		.out_col (out_col_13_17),
		.out_data (out_data_13_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_18;
	wire signed [DATA_WIDTH-1:0] out_col_13_18;
	wire signed [DATA_WIDTH-1:0] out_data_13_18;
	integer_mac_pe mac_pe_13_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_17),
		.in_col (out_col_12_18),
		.out_row (out_row_13_18),
		.out_col (out_col_13_18),
		.out_data (out_data_13_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_19;
	wire signed [DATA_WIDTH-1:0] out_col_13_19;
	wire signed [DATA_WIDTH-1:0] out_data_13_19;
	integer_mac_pe mac_pe_13_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_18),
		.in_col (out_col_12_19),
		.out_row (out_row_13_19),
		.out_col (out_col_13_19),
		.out_data (out_data_13_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_20;
	wire signed [DATA_WIDTH-1:0] out_col_13_20;
	wire signed [DATA_WIDTH-1:0] out_data_13_20;
	integer_mac_pe mac_pe_13_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_19),
		.in_col (out_col_12_20),
		.out_row (out_row_13_20),
		.out_col (out_col_13_20),
		.out_data (out_data_13_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_21;
	wire signed [DATA_WIDTH-1:0] out_col_13_21;
	wire signed [DATA_WIDTH-1:0] out_data_13_21;
	integer_mac_pe mac_pe_13_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_20),
		.in_col (out_col_12_21),
		.out_row (out_row_13_21),
		.out_col (out_col_13_21),
		.out_data (out_data_13_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_22;
	wire signed [DATA_WIDTH-1:0] out_col_13_22;
	wire signed [DATA_WIDTH-1:0] out_data_13_22;
	integer_mac_pe mac_pe_13_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_21),
		.in_col (out_col_12_22),
		.out_row (out_row_13_22),
		.out_col (out_col_13_22),
		.out_data (out_data_13_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_23;
	wire signed [DATA_WIDTH-1:0] out_col_13_23;
	wire signed [DATA_WIDTH-1:0] out_data_13_23;
	integer_mac_pe mac_pe_13_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_22),
		.in_col (out_col_12_23),
		.out_row (out_row_13_23),
		.out_col (out_col_13_23),
		.out_data (out_data_13_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_24;
	wire signed [DATA_WIDTH-1:0] out_col_13_24;
	wire signed [DATA_WIDTH-1:0] out_data_13_24;
	integer_mac_pe mac_pe_13_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_23),
		.in_col (out_col_12_24),
		.out_row (out_row_13_24),
		.out_col (out_col_13_24),
		.out_data (out_data_13_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_25;
	wire signed [DATA_WIDTH-1:0] out_col_13_25;
	wire signed [DATA_WIDTH-1:0] out_data_13_25;
	integer_mac_pe mac_pe_13_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_24),
		.in_col (out_col_12_25),
		.out_row (out_row_13_25),
		.out_col (out_col_13_25),
		.out_data (out_data_13_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_26;
	wire signed [DATA_WIDTH-1:0] out_col_13_26;
	wire signed [DATA_WIDTH-1:0] out_data_13_26;
	integer_mac_pe mac_pe_13_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_25),
		.in_col (out_col_12_26),
		.out_row (out_row_13_26),
		.out_col (out_col_13_26),
		.out_data (out_data_13_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_27;
	wire signed [DATA_WIDTH-1:0] out_col_13_27;
	wire signed [DATA_WIDTH-1:0] out_data_13_27;
	integer_mac_pe mac_pe_13_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_26),
		.in_col (out_col_12_27),
		.out_row (out_row_13_27),
		.out_col (out_col_13_27),
		.out_data (out_data_13_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_28;
	wire signed [DATA_WIDTH-1:0] out_col_13_28;
	wire signed [DATA_WIDTH-1:0] out_data_13_28;
	integer_mac_pe mac_pe_13_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_27),
		.in_col (out_col_12_28),
		.out_row (out_row_13_28),
		.out_col (out_col_13_28),
		.out_data (out_data_13_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_29;
	wire signed [DATA_WIDTH-1:0] out_col_13_29;
	wire signed [DATA_WIDTH-1:0] out_data_13_29;
	integer_mac_pe mac_pe_13_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_28),
		.in_col (out_col_12_29),
		.out_row (out_row_13_29),
		.out_col (out_col_13_29),
		.out_data (out_data_13_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_30;
	wire signed [DATA_WIDTH-1:0] out_col_13_30;
	wire signed [DATA_WIDTH-1:0] out_data_13_30;
	integer_mac_pe mac_pe_13_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_29),
		.in_col (out_col_12_30),
		.out_row (out_row_13_30),
		.out_col (out_col_13_30),
		.out_data (out_data_13_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_13_31;
	wire signed [DATA_WIDTH-1:0] out_col_13_31;
	wire signed [DATA_WIDTH-1:0] out_data_13_31;
	integer_mac_pe mac_pe_13_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_13_30),
		.in_col (out_col_12_31),
		.out_row (out_row_13_31),
		.out_col (out_col_13_31),
		.out_data (out_data_13_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_0;
	wire signed [DATA_WIDTH-1:0] out_col_14_0;
	wire signed [DATA_WIDTH-1:0] out_data_14_0;
	integer_mac_pe mac_pe_14_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_14_out),
		.in_col (out_col_13_0),
		.out_row (out_row_14_0),
		.out_col (out_col_14_0),
		.out_data (out_data_14_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_1;
	wire signed [DATA_WIDTH-1:0] out_col_14_1;
	wire signed [DATA_WIDTH-1:0] out_data_14_1;
	integer_mac_pe mac_pe_14_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_0),
		.in_col (out_col_13_1),
		.out_row (out_row_14_1),
		.out_col (out_col_14_1),
		.out_data (out_data_14_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_2;
	wire signed [DATA_WIDTH-1:0] out_col_14_2;
	wire signed [DATA_WIDTH-1:0] out_data_14_2;
	integer_mac_pe mac_pe_14_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_1),
		.in_col (out_col_13_2),
		.out_row (out_row_14_2),
		.out_col (out_col_14_2),
		.out_data (out_data_14_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_3;
	wire signed [DATA_WIDTH-1:0] out_col_14_3;
	wire signed [DATA_WIDTH-1:0] out_data_14_3;
	integer_mac_pe mac_pe_14_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_2),
		.in_col (out_col_13_3),
		.out_row (out_row_14_3),
		.out_col (out_col_14_3),
		.out_data (out_data_14_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_4;
	wire signed [DATA_WIDTH-1:0] out_col_14_4;
	wire signed [DATA_WIDTH-1:0] out_data_14_4;
	integer_mac_pe mac_pe_14_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_3),
		.in_col (out_col_13_4),
		.out_row (out_row_14_4),
		.out_col (out_col_14_4),
		.out_data (out_data_14_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_5;
	wire signed [DATA_WIDTH-1:0] out_col_14_5;
	wire signed [DATA_WIDTH-1:0] out_data_14_5;
	integer_mac_pe mac_pe_14_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_4),
		.in_col (out_col_13_5),
		.out_row (out_row_14_5),
		.out_col (out_col_14_5),
		.out_data (out_data_14_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_6;
	wire signed [DATA_WIDTH-1:0] out_col_14_6;
	wire signed [DATA_WIDTH-1:0] out_data_14_6;
	integer_mac_pe mac_pe_14_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_5),
		.in_col (out_col_13_6),
		.out_row (out_row_14_6),
		.out_col (out_col_14_6),
		.out_data (out_data_14_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_7;
	wire signed [DATA_WIDTH-1:0] out_col_14_7;
	wire signed [DATA_WIDTH-1:0] out_data_14_7;
	integer_mac_pe mac_pe_14_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_6),
		.in_col (out_col_13_7),
		.out_row (out_row_14_7),
		.out_col (out_col_14_7),
		.out_data (out_data_14_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_8;
	wire signed [DATA_WIDTH-1:0] out_col_14_8;
	wire signed [DATA_WIDTH-1:0] out_data_14_8;
	integer_mac_pe mac_pe_14_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_7),
		.in_col (out_col_13_8),
		.out_row (out_row_14_8),
		.out_col (out_col_14_8),
		.out_data (out_data_14_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_9;
	wire signed [DATA_WIDTH-1:0] out_col_14_9;
	wire signed [DATA_WIDTH-1:0] out_data_14_9;
	integer_mac_pe mac_pe_14_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_8),
		.in_col (out_col_13_9),
		.out_row (out_row_14_9),
		.out_col (out_col_14_9),
		.out_data (out_data_14_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_10;
	wire signed [DATA_WIDTH-1:0] out_col_14_10;
	wire signed [DATA_WIDTH-1:0] out_data_14_10;
	integer_mac_pe mac_pe_14_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_9),
		.in_col (out_col_13_10),
		.out_row (out_row_14_10),
		.out_col (out_col_14_10),
		.out_data (out_data_14_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_11;
	wire signed [DATA_WIDTH-1:0] out_col_14_11;
	wire signed [DATA_WIDTH-1:0] out_data_14_11;
	integer_mac_pe mac_pe_14_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_10),
		.in_col (out_col_13_11),
		.out_row (out_row_14_11),
		.out_col (out_col_14_11),
		.out_data (out_data_14_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_12;
	wire signed [DATA_WIDTH-1:0] out_col_14_12;
	wire signed [DATA_WIDTH-1:0] out_data_14_12;
	integer_mac_pe mac_pe_14_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_11),
		.in_col (out_col_13_12),
		.out_row (out_row_14_12),
		.out_col (out_col_14_12),
		.out_data (out_data_14_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_13;
	wire signed [DATA_WIDTH-1:0] out_col_14_13;
	wire signed [DATA_WIDTH-1:0] out_data_14_13;
	integer_mac_pe mac_pe_14_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_12),
		.in_col (out_col_13_13),
		.out_row (out_row_14_13),
		.out_col (out_col_14_13),
		.out_data (out_data_14_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_14;
	wire signed [DATA_WIDTH-1:0] out_col_14_14;
	wire signed [DATA_WIDTH-1:0] out_data_14_14;
	integer_mac_pe mac_pe_14_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_13),
		.in_col (out_col_13_14),
		.out_row (out_row_14_14),
		.out_col (out_col_14_14),
		.out_data (out_data_14_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_15;
	wire signed [DATA_WIDTH-1:0] out_col_14_15;
	wire signed [DATA_WIDTH-1:0] out_data_14_15;
	integer_mac_pe mac_pe_14_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_14),
		.in_col (out_col_13_15),
		.out_row (out_row_14_15),
		.out_col (out_col_14_15),
		.out_data (out_data_14_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_16;
	wire signed [DATA_WIDTH-1:0] out_col_14_16;
	wire signed [DATA_WIDTH-1:0] out_data_14_16;
	integer_mac_pe mac_pe_14_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_15),
		.in_col (out_col_13_16),
		.out_row (out_row_14_16),
		.out_col (out_col_14_16),
		.out_data (out_data_14_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_17;
	wire signed [DATA_WIDTH-1:0] out_col_14_17;
	wire signed [DATA_WIDTH-1:0] out_data_14_17;
	integer_mac_pe mac_pe_14_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_16),
		.in_col (out_col_13_17),
		.out_row (out_row_14_17),
		.out_col (out_col_14_17),
		.out_data (out_data_14_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_18;
	wire signed [DATA_WIDTH-1:0] out_col_14_18;
	wire signed [DATA_WIDTH-1:0] out_data_14_18;
	integer_mac_pe mac_pe_14_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_17),
		.in_col (out_col_13_18),
		.out_row (out_row_14_18),
		.out_col (out_col_14_18),
		.out_data (out_data_14_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_19;
	wire signed [DATA_WIDTH-1:0] out_col_14_19;
	wire signed [DATA_WIDTH-1:0] out_data_14_19;
	integer_mac_pe mac_pe_14_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_18),
		.in_col (out_col_13_19),
		.out_row (out_row_14_19),
		.out_col (out_col_14_19),
		.out_data (out_data_14_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_20;
	wire signed [DATA_WIDTH-1:0] out_col_14_20;
	wire signed [DATA_WIDTH-1:0] out_data_14_20;
	integer_mac_pe mac_pe_14_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_19),
		.in_col (out_col_13_20),
		.out_row (out_row_14_20),
		.out_col (out_col_14_20),
		.out_data (out_data_14_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_21;
	wire signed [DATA_WIDTH-1:0] out_col_14_21;
	wire signed [DATA_WIDTH-1:0] out_data_14_21;
	integer_mac_pe mac_pe_14_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_20),
		.in_col (out_col_13_21),
		.out_row (out_row_14_21),
		.out_col (out_col_14_21),
		.out_data (out_data_14_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_22;
	wire signed [DATA_WIDTH-1:0] out_col_14_22;
	wire signed [DATA_WIDTH-1:0] out_data_14_22;
	integer_mac_pe mac_pe_14_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_21),
		.in_col (out_col_13_22),
		.out_row (out_row_14_22),
		.out_col (out_col_14_22),
		.out_data (out_data_14_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_23;
	wire signed [DATA_WIDTH-1:0] out_col_14_23;
	wire signed [DATA_WIDTH-1:0] out_data_14_23;
	integer_mac_pe mac_pe_14_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_22),
		.in_col (out_col_13_23),
		.out_row (out_row_14_23),
		.out_col (out_col_14_23),
		.out_data (out_data_14_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_24;
	wire signed [DATA_WIDTH-1:0] out_col_14_24;
	wire signed [DATA_WIDTH-1:0] out_data_14_24;
	integer_mac_pe mac_pe_14_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_23),
		.in_col (out_col_13_24),
		.out_row (out_row_14_24),
		.out_col (out_col_14_24),
		.out_data (out_data_14_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_25;
	wire signed [DATA_WIDTH-1:0] out_col_14_25;
	wire signed [DATA_WIDTH-1:0] out_data_14_25;
	integer_mac_pe mac_pe_14_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_24),
		.in_col (out_col_13_25),
		.out_row (out_row_14_25),
		.out_col (out_col_14_25),
		.out_data (out_data_14_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_26;
	wire signed [DATA_WIDTH-1:0] out_col_14_26;
	wire signed [DATA_WIDTH-1:0] out_data_14_26;
	integer_mac_pe mac_pe_14_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_25),
		.in_col (out_col_13_26),
		.out_row (out_row_14_26),
		.out_col (out_col_14_26),
		.out_data (out_data_14_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_27;
	wire signed [DATA_WIDTH-1:0] out_col_14_27;
	wire signed [DATA_WIDTH-1:0] out_data_14_27;
	integer_mac_pe mac_pe_14_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_26),
		.in_col (out_col_13_27),
		.out_row (out_row_14_27),
		.out_col (out_col_14_27),
		.out_data (out_data_14_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_28;
	wire signed [DATA_WIDTH-1:0] out_col_14_28;
	wire signed [DATA_WIDTH-1:0] out_data_14_28;
	integer_mac_pe mac_pe_14_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_27),
		.in_col (out_col_13_28),
		.out_row (out_row_14_28),
		.out_col (out_col_14_28),
		.out_data (out_data_14_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_29;
	wire signed [DATA_WIDTH-1:0] out_col_14_29;
	wire signed [DATA_WIDTH-1:0] out_data_14_29;
	integer_mac_pe mac_pe_14_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_28),
		.in_col (out_col_13_29),
		.out_row (out_row_14_29),
		.out_col (out_col_14_29),
		.out_data (out_data_14_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_30;
	wire signed [DATA_WIDTH-1:0] out_col_14_30;
	wire signed [DATA_WIDTH-1:0] out_data_14_30;
	integer_mac_pe mac_pe_14_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_29),
		.in_col (out_col_13_30),
		.out_row (out_row_14_30),
		.out_col (out_col_14_30),
		.out_data (out_data_14_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_14_31;
	wire signed [DATA_WIDTH-1:0] out_col_14_31;
	wire signed [DATA_WIDTH-1:0] out_data_14_31;
	integer_mac_pe mac_pe_14_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_14_30),
		.in_col (out_col_13_31),
		.out_row (out_row_14_31),
		.out_col (out_col_14_31),
		.out_data (out_data_14_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_0;
	wire signed [DATA_WIDTH-1:0] out_col_15_0;
	wire signed [DATA_WIDTH-1:0] out_data_15_0;
	integer_mac_pe mac_pe_15_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_15_out),
		.in_col (out_col_14_0),
		.out_row (out_row_15_0),
		.out_col (out_col_15_0),
		.out_data (out_data_15_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_1;
	wire signed [DATA_WIDTH-1:0] out_col_15_1;
	wire signed [DATA_WIDTH-1:0] out_data_15_1;
	integer_mac_pe mac_pe_15_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_0),
		.in_col (out_col_14_1),
		.out_row (out_row_15_1),
		.out_col (out_col_15_1),
		.out_data (out_data_15_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_2;
	wire signed [DATA_WIDTH-1:0] out_col_15_2;
	wire signed [DATA_WIDTH-1:0] out_data_15_2;
	integer_mac_pe mac_pe_15_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_1),
		.in_col (out_col_14_2),
		.out_row (out_row_15_2),
		.out_col (out_col_15_2),
		.out_data (out_data_15_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_3;
	wire signed [DATA_WIDTH-1:0] out_col_15_3;
	wire signed [DATA_WIDTH-1:0] out_data_15_3;
	integer_mac_pe mac_pe_15_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_2),
		.in_col (out_col_14_3),
		.out_row (out_row_15_3),
		.out_col (out_col_15_3),
		.out_data (out_data_15_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_4;
	wire signed [DATA_WIDTH-1:0] out_col_15_4;
	wire signed [DATA_WIDTH-1:0] out_data_15_4;
	integer_mac_pe mac_pe_15_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_3),
		.in_col (out_col_14_4),
		.out_row (out_row_15_4),
		.out_col (out_col_15_4),
		.out_data (out_data_15_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_5;
	wire signed [DATA_WIDTH-1:0] out_col_15_5;
	wire signed [DATA_WIDTH-1:0] out_data_15_5;
	integer_mac_pe mac_pe_15_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_4),
		.in_col (out_col_14_5),
		.out_row (out_row_15_5),
		.out_col (out_col_15_5),
		.out_data (out_data_15_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_6;
	wire signed [DATA_WIDTH-1:0] out_col_15_6;
	wire signed [DATA_WIDTH-1:0] out_data_15_6;
	integer_mac_pe mac_pe_15_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_5),
		.in_col (out_col_14_6),
		.out_row (out_row_15_6),
		.out_col (out_col_15_6),
		.out_data (out_data_15_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_7;
	wire signed [DATA_WIDTH-1:0] out_col_15_7;
	wire signed [DATA_WIDTH-1:0] out_data_15_7;
	integer_mac_pe mac_pe_15_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_6),
		.in_col (out_col_14_7),
		.out_row (out_row_15_7),
		.out_col (out_col_15_7),
		.out_data (out_data_15_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_8;
	wire signed [DATA_WIDTH-1:0] out_col_15_8;
	wire signed [DATA_WIDTH-1:0] out_data_15_8;
	integer_mac_pe mac_pe_15_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_7),
		.in_col (out_col_14_8),
		.out_row (out_row_15_8),
		.out_col (out_col_15_8),
		.out_data (out_data_15_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_9;
	wire signed [DATA_WIDTH-1:0] out_col_15_9;
	wire signed [DATA_WIDTH-1:0] out_data_15_9;
	integer_mac_pe mac_pe_15_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_8),
		.in_col (out_col_14_9),
		.out_row (out_row_15_9),
		.out_col (out_col_15_9),
		.out_data (out_data_15_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_10;
	wire signed [DATA_WIDTH-1:0] out_col_15_10;
	wire signed [DATA_WIDTH-1:0] out_data_15_10;
	integer_mac_pe mac_pe_15_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_9),
		.in_col (out_col_14_10),
		.out_row (out_row_15_10),
		.out_col (out_col_15_10),
		.out_data (out_data_15_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_11;
	wire signed [DATA_WIDTH-1:0] out_col_15_11;
	wire signed [DATA_WIDTH-1:0] out_data_15_11;
	integer_mac_pe mac_pe_15_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_10),
		.in_col (out_col_14_11),
		.out_row (out_row_15_11),
		.out_col (out_col_15_11),
		.out_data (out_data_15_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_12;
	wire signed [DATA_WIDTH-1:0] out_col_15_12;
	wire signed [DATA_WIDTH-1:0] out_data_15_12;
	integer_mac_pe mac_pe_15_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_11),
		.in_col (out_col_14_12),
		.out_row (out_row_15_12),
		.out_col (out_col_15_12),
		.out_data (out_data_15_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_13;
	wire signed [DATA_WIDTH-1:0] out_col_15_13;
	wire signed [DATA_WIDTH-1:0] out_data_15_13;
	integer_mac_pe mac_pe_15_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_12),
		.in_col (out_col_14_13),
		.out_row (out_row_15_13),
		.out_col (out_col_15_13),
		.out_data (out_data_15_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_14;
	wire signed [DATA_WIDTH-1:0] out_col_15_14;
	wire signed [DATA_WIDTH-1:0] out_data_15_14;
	integer_mac_pe mac_pe_15_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_13),
		.in_col (out_col_14_14),
		.out_row (out_row_15_14),
		.out_col (out_col_15_14),
		.out_data (out_data_15_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_15;
	wire signed [DATA_WIDTH-1:0] out_col_15_15;
	wire signed [DATA_WIDTH-1:0] out_data_15_15;
	integer_mac_pe mac_pe_15_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_14),
		.in_col (out_col_14_15),
		.out_row (out_row_15_15),
		.out_col (out_col_15_15),
		.out_data (out_data_15_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_16;
	wire signed [DATA_WIDTH-1:0] out_col_15_16;
	wire signed [DATA_WIDTH-1:0] out_data_15_16;
	integer_mac_pe mac_pe_15_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_15),
		.in_col (out_col_14_16),
		.out_row (out_row_15_16),
		.out_col (out_col_15_16),
		.out_data (out_data_15_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_17;
	wire signed [DATA_WIDTH-1:0] out_col_15_17;
	wire signed [DATA_WIDTH-1:0] out_data_15_17;
	integer_mac_pe mac_pe_15_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_16),
		.in_col (out_col_14_17),
		.out_row (out_row_15_17),
		.out_col (out_col_15_17),
		.out_data (out_data_15_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_18;
	wire signed [DATA_WIDTH-1:0] out_col_15_18;
	wire signed [DATA_WIDTH-1:0] out_data_15_18;
	integer_mac_pe mac_pe_15_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_17),
		.in_col (out_col_14_18),
		.out_row (out_row_15_18),
		.out_col (out_col_15_18),
		.out_data (out_data_15_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_19;
	wire signed [DATA_WIDTH-1:0] out_col_15_19;
	wire signed [DATA_WIDTH-1:0] out_data_15_19;
	integer_mac_pe mac_pe_15_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_18),
		.in_col (out_col_14_19),
		.out_row (out_row_15_19),
		.out_col (out_col_15_19),
		.out_data (out_data_15_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_20;
	wire signed [DATA_WIDTH-1:0] out_col_15_20;
	wire signed [DATA_WIDTH-1:0] out_data_15_20;
	integer_mac_pe mac_pe_15_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_19),
		.in_col (out_col_14_20),
		.out_row (out_row_15_20),
		.out_col (out_col_15_20),
		.out_data (out_data_15_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_21;
	wire signed [DATA_WIDTH-1:0] out_col_15_21;
	wire signed [DATA_WIDTH-1:0] out_data_15_21;
	integer_mac_pe mac_pe_15_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_20),
		.in_col (out_col_14_21),
		.out_row (out_row_15_21),
		.out_col (out_col_15_21),
		.out_data (out_data_15_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_22;
	wire signed [DATA_WIDTH-1:0] out_col_15_22;
	wire signed [DATA_WIDTH-1:0] out_data_15_22;
	integer_mac_pe mac_pe_15_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_21),
		.in_col (out_col_14_22),
		.out_row (out_row_15_22),
		.out_col (out_col_15_22),
		.out_data (out_data_15_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_23;
	wire signed [DATA_WIDTH-1:0] out_col_15_23;
	wire signed [DATA_WIDTH-1:0] out_data_15_23;
	integer_mac_pe mac_pe_15_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_22),
		.in_col (out_col_14_23),
		.out_row (out_row_15_23),
		.out_col (out_col_15_23),
		.out_data (out_data_15_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_24;
	wire signed [DATA_WIDTH-1:0] out_col_15_24;
	wire signed [DATA_WIDTH-1:0] out_data_15_24;
	integer_mac_pe mac_pe_15_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_23),
		.in_col (out_col_14_24),
		.out_row (out_row_15_24),
		.out_col (out_col_15_24),
		.out_data (out_data_15_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_25;
	wire signed [DATA_WIDTH-1:0] out_col_15_25;
	wire signed [DATA_WIDTH-1:0] out_data_15_25;
	integer_mac_pe mac_pe_15_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_24),
		.in_col (out_col_14_25),
		.out_row (out_row_15_25),
		.out_col (out_col_15_25),
		.out_data (out_data_15_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_26;
	wire signed [DATA_WIDTH-1:0] out_col_15_26;
	wire signed [DATA_WIDTH-1:0] out_data_15_26;
	integer_mac_pe mac_pe_15_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_25),
		.in_col (out_col_14_26),
		.out_row (out_row_15_26),
		.out_col (out_col_15_26),
		.out_data (out_data_15_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_27;
	wire signed [DATA_WIDTH-1:0] out_col_15_27;
	wire signed [DATA_WIDTH-1:0] out_data_15_27;
	integer_mac_pe mac_pe_15_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_26),
		.in_col (out_col_14_27),
		.out_row (out_row_15_27),
		.out_col (out_col_15_27),
		.out_data (out_data_15_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_28;
	wire signed [DATA_WIDTH-1:0] out_col_15_28;
	wire signed [DATA_WIDTH-1:0] out_data_15_28;
	integer_mac_pe mac_pe_15_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_27),
		.in_col (out_col_14_28),
		.out_row (out_row_15_28),
		.out_col (out_col_15_28),
		.out_data (out_data_15_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_29;
	wire signed [DATA_WIDTH-1:0] out_col_15_29;
	wire signed [DATA_WIDTH-1:0] out_data_15_29;
	integer_mac_pe mac_pe_15_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_28),
		.in_col (out_col_14_29),
		.out_row (out_row_15_29),
		.out_col (out_col_15_29),
		.out_data (out_data_15_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_30;
	wire signed [DATA_WIDTH-1:0] out_col_15_30;
	wire signed [DATA_WIDTH-1:0] out_data_15_30;
	integer_mac_pe mac_pe_15_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_29),
		.in_col (out_col_14_30),
		.out_row (out_row_15_30),
		.out_col (out_col_15_30),
		.out_data (out_data_15_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_15_31;
	wire signed [DATA_WIDTH-1:0] out_col_15_31;
	wire signed [DATA_WIDTH-1:0] out_data_15_31;
	integer_mac_pe mac_pe_15_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_15_30),
		.in_col (out_col_14_31),
		.out_row (out_row_15_31),
		.out_col (out_col_15_31),
		.out_data (out_data_15_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_0;
	wire signed [DATA_WIDTH-1:0] out_col_16_0;
	wire signed [DATA_WIDTH-1:0] out_data_16_0;
	integer_mac_pe mac_pe_16_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_16_out),
		.in_col (out_col_15_0),
		.out_row (out_row_16_0),
		.out_col (out_col_16_0),
		.out_data (out_data_16_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_1;
	wire signed [DATA_WIDTH-1:0] out_col_16_1;
	wire signed [DATA_WIDTH-1:0] out_data_16_1;
	integer_mac_pe mac_pe_16_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_0),
		.in_col (out_col_15_1),
		.out_row (out_row_16_1),
		.out_col (out_col_16_1),
		.out_data (out_data_16_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_2;
	wire signed [DATA_WIDTH-1:0] out_col_16_2;
	wire signed [DATA_WIDTH-1:0] out_data_16_2;
	integer_mac_pe mac_pe_16_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_1),
		.in_col (out_col_15_2),
		.out_row (out_row_16_2),
		.out_col (out_col_16_2),
		.out_data (out_data_16_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_3;
	wire signed [DATA_WIDTH-1:0] out_col_16_3;
	wire signed [DATA_WIDTH-1:0] out_data_16_3;
	integer_mac_pe mac_pe_16_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_2),
		.in_col (out_col_15_3),
		.out_row (out_row_16_3),
		.out_col (out_col_16_3),
		.out_data (out_data_16_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_4;
	wire signed [DATA_WIDTH-1:0] out_col_16_4;
	wire signed [DATA_WIDTH-1:0] out_data_16_4;
	integer_mac_pe mac_pe_16_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_3),
		.in_col (out_col_15_4),
		.out_row (out_row_16_4),
		.out_col (out_col_16_4),
		.out_data (out_data_16_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_5;
	wire signed [DATA_WIDTH-1:0] out_col_16_5;
	wire signed [DATA_WIDTH-1:0] out_data_16_5;
	integer_mac_pe mac_pe_16_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_4),
		.in_col (out_col_15_5),
		.out_row (out_row_16_5),
		.out_col (out_col_16_5),
		.out_data (out_data_16_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_6;
	wire signed [DATA_WIDTH-1:0] out_col_16_6;
	wire signed [DATA_WIDTH-1:0] out_data_16_6;
	integer_mac_pe mac_pe_16_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_5),
		.in_col (out_col_15_6),
		.out_row (out_row_16_6),
		.out_col (out_col_16_6),
		.out_data (out_data_16_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_7;
	wire signed [DATA_WIDTH-1:0] out_col_16_7;
	wire signed [DATA_WIDTH-1:0] out_data_16_7;
	integer_mac_pe mac_pe_16_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_6),
		.in_col (out_col_15_7),
		.out_row (out_row_16_7),
		.out_col (out_col_16_7),
		.out_data (out_data_16_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_8;
	wire signed [DATA_WIDTH-1:0] out_col_16_8;
	wire signed [DATA_WIDTH-1:0] out_data_16_8;
	integer_mac_pe mac_pe_16_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_7),
		.in_col (out_col_15_8),
		.out_row (out_row_16_8),
		.out_col (out_col_16_8),
		.out_data (out_data_16_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_9;
	wire signed [DATA_WIDTH-1:0] out_col_16_9;
	wire signed [DATA_WIDTH-1:0] out_data_16_9;
	integer_mac_pe mac_pe_16_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_8),
		.in_col (out_col_15_9),
		.out_row (out_row_16_9),
		.out_col (out_col_16_9),
		.out_data (out_data_16_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_10;
	wire signed [DATA_WIDTH-1:0] out_col_16_10;
	wire signed [DATA_WIDTH-1:0] out_data_16_10;
	integer_mac_pe mac_pe_16_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_9),
		.in_col (out_col_15_10),
		.out_row (out_row_16_10),
		.out_col (out_col_16_10),
		.out_data (out_data_16_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_11;
	wire signed [DATA_WIDTH-1:0] out_col_16_11;
	wire signed [DATA_WIDTH-1:0] out_data_16_11;
	integer_mac_pe mac_pe_16_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_10),
		.in_col (out_col_15_11),
		.out_row (out_row_16_11),
		.out_col (out_col_16_11),
		.out_data (out_data_16_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_12;
	wire signed [DATA_WIDTH-1:0] out_col_16_12;
	wire signed [DATA_WIDTH-1:0] out_data_16_12;
	integer_mac_pe mac_pe_16_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_11),
		.in_col (out_col_15_12),
		.out_row (out_row_16_12),
		.out_col (out_col_16_12),
		.out_data (out_data_16_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_13;
	wire signed [DATA_WIDTH-1:0] out_col_16_13;
	wire signed [DATA_WIDTH-1:0] out_data_16_13;
	integer_mac_pe mac_pe_16_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_12),
		.in_col (out_col_15_13),
		.out_row (out_row_16_13),
		.out_col (out_col_16_13),
		.out_data (out_data_16_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_14;
	wire signed [DATA_WIDTH-1:0] out_col_16_14;
	wire signed [DATA_WIDTH-1:0] out_data_16_14;
	integer_mac_pe mac_pe_16_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_13),
		.in_col (out_col_15_14),
		.out_row (out_row_16_14),
		.out_col (out_col_16_14),
		.out_data (out_data_16_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_15;
	wire signed [DATA_WIDTH-1:0] out_col_16_15;
	wire signed [DATA_WIDTH-1:0] out_data_16_15;
	integer_mac_pe mac_pe_16_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_14),
		.in_col (out_col_15_15),
		.out_row (out_row_16_15),
		.out_col (out_col_16_15),
		.out_data (out_data_16_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_16;
	wire signed [DATA_WIDTH-1:0] out_col_16_16;
	wire signed [DATA_WIDTH-1:0] out_data_16_16;
	integer_mac_pe mac_pe_16_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_15),
		.in_col (out_col_15_16),
		.out_row (out_row_16_16),
		.out_col (out_col_16_16),
		.out_data (out_data_16_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_17;
	wire signed [DATA_WIDTH-1:0] out_col_16_17;
	wire signed [DATA_WIDTH-1:0] out_data_16_17;
	integer_mac_pe mac_pe_16_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_16),
		.in_col (out_col_15_17),
		.out_row (out_row_16_17),
		.out_col (out_col_16_17),
		.out_data (out_data_16_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_18;
	wire signed [DATA_WIDTH-1:0] out_col_16_18;
	wire signed [DATA_WIDTH-1:0] out_data_16_18;
	integer_mac_pe mac_pe_16_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_17),
		.in_col (out_col_15_18),
		.out_row (out_row_16_18),
		.out_col (out_col_16_18),
		.out_data (out_data_16_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_19;
	wire signed [DATA_WIDTH-1:0] out_col_16_19;
	wire signed [DATA_WIDTH-1:0] out_data_16_19;
	integer_mac_pe mac_pe_16_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_18),
		.in_col (out_col_15_19),
		.out_row (out_row_16_19),
		.out_col (out_col_16_19),
		.out_data (out_data_16_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_20;
	wire signed [DATA_WIDTH-1:0] out_col_16_20;
	wire signed [DATA_WIDTH-1:0] out_data_16_20;
	integer_mac_pe mac_pe_16_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_19),
		.in_col (out_col_15_20),
		.out_row (out_row_16_20),
		.out_col (out_col_16_20),
		.out_data (out_data_16_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_21;
	wire signed [DATA_WIDTH-1:0] out_col_16_21;
	wire signed [DATA_WIDTH-1:0] out_data_16_21;
	integer_mac_pe mac_pe_16_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_20),
		.in_col (out_col_15_21),
		.out_row (out_row_16_21),
		.out_col (out_col_16_21),
		.out_data (out_data_16_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_22;
	wire signed [DATA_WIDTH-1:0] out_col_16_22;
	wire signed [DATA_WIDTH-1:0] out_data_16_22;
	integer_mac_pe mac_pe_16_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_21),
		.in_col (out_col_15_22),
		.out_row (out_row_16_22),
		.out_col (out_col_16_22),
		.out_data (out_data_16_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_23;
	wire signed [DATA_WIDTH-1:0] out_col_16_23;
	wire signed [DATA_WIDTH-1:0] out_data_16_23;
	integer_mac_pe mac_pe_16_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_22),
		.in_col (out_col_15_23),
		.out_row (out_row_16_23),
		.out_col (out_col_16_23),
		.out_data (out_data_16_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_24;
	wire signed [DATA_WIDTH-1:0] out_col_16_24;
	wire signed [DATA_WIDTH-1:0] out_data_16_24;
	integer_mac_pe mac_pe_16_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_23),
		.in_col (out_col_15_24),
		.out_row (out_row_16_24),
		.out_col (out_col_16_24),
		.out_data (out_data_16_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_25;
	wire signed [DATA_WIDTH-1:0] out_col_16_25;
	wire signed [DATA_WIDTH-1:0] out_data_16_25;
	integer_mac_pe mac_pe_16_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_24),
		.in_col (out_col_15_25),
		.out_row (out_row_16_25),
		.out_col (out_col_16_25),
		.out_data (out_data_16_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_26;
	wire signed [DATA_WIDTH-1:0] out_col_16_26;
	wire signed [DATA_WIDTH-1:0] out_data_16_26;
	integer_mac_pe mac_pe_16_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_25),
		.in_col (out_col_15_26),
		.out_row (out_row_16_26),
		.out_col (out_col_16_26),
		.out_data (out_data_16_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_27;
	wire signed [DATA_WIDTH-1:0] out_col_16_27;
	wire signed [DATA_WIDTH-1:0] out_data_16_27;
	integer_mac_pe mac_pe_16_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_26),
		.in_col (out_col_15_27),
		.out_row (out_row_16_27),
		.out_col (out_col_16_27),
		.out_data (out_data_16_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_28;
	wire signed [DATA_WIDTH-1:0] out_col_16_28;
	wire signed [DATA_WIDTH-1:0] out_data_16_28;
	integer_mac_pe mac_pe_16_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_27),
		.in_col (out_col_15_28),
		.out_row (out_row_16_28),
		.out_col (out_col_16_28),
		.out_data (out_data_16_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_29;
	wire signed [DATA_WIDTH-1:0] out_col_16_29;
	wire signed [DATA_WIDTH-1:0] out_data_16_29;
	integer_mac_pe mac_pe_16_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_28),
		.in_col (out_col_15_29),
		.out_row (out_row_16_29),
		.out_col (out_col_16_29),
		.out_data (out_data_16_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_30;
	wire signed [DATA_WIDTH-1:0] out_col_16_30;
	wire signed [DATA_WIDTH-1:0] out_data_16_30;
	integer_mac_pe mac_pe_16_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_29),
		.in_col (out_col_15_30),
		.out_row (out_row_16_30),
		.out_col (out_col_16_30),
		.out_data (out_data_16_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_16_31;
	wire signed [DATA_WIDTH-1:0] out_col_16_31;
	wire signed [DATA_WIDTH-1:0] out_data_16_31;
	integer_mac_pe mac_pe_16_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_16_30),
		.in_col (out_col_15_31),
		.out_row (out_row_16_31),
		.out_col (out_col_16_31),
		.out_data (out_data_16_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_0;
	wire signed [DATA_WIDTH-1:0] out_col_17_0;
	wire signed [DATA_WIDTH-1:0] out_data_17_0;
	integer_mac_pe mac_pe_17_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_17_out),
		.in_col (out_col_16_0),
		.out_row (out_row_17_0),
		.out_col (out_col_17_0),
		.out_data (out_data_17_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_1;
	wire signed [DATA_WIDTH-1:0] out_col_17_1;
	wire signed [DATA_WIDTH-1:0] out_data_17_1;
	integer_mac_pe mac_pe_17_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_0),
		.in_col (out_col_16_1),
		.out_row (out_row_17_1),
		.out_col (out_col_17_1),
		.out_data (out_data_17_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_2;
	wire signed [DATA_WIDTH-1:0] out_col_17_2;
	wire signed [DATA_WIDTH-1:0] out_data_17_2;
	integer_mac_pe mac_pe_17_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_1),
		.in_col (out_col_16_2),
		.out_row (out_row_17_2),
		.out_col (out_col_17_2),
		.out_data (out_data_17_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_3;
	wire signed [DATA_WIDTH-1:0] out_col_17_3;
	wire signed [DATA_WIDTH-1:0] out_data_17_3;
	integer_mac_pe mac_pe_17_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_2),
		.in_col (out_col_16_3),
		.out_row (out_row_17_3),
		.out_col (out_col_17_3),
		.out_data (out_data_17_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_4;
	wire signed [DATA_WIDTH-1:0] out_col_17_4;
	wire signed [DATA_WIDTH-1:0] out_data_17_4;
	integer_mac_pe mac_pe_17_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_3),
		.in_col (out_col_16_4),
		.out_row (out_row_17_4),
		.out_col (out_col_17_4),
		.out_data (out_data_17_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_5;
	wire signed [DATA_WIDTH-1:0] out_col_17_5;
	wire signed [DATA_WIDTH-1:0] out_data_17_5;
	integer_mac_pe mac_pe_17_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_4),
		.in_col (out_col_16_5),
		.out_row (out_row_17_5),
		.out_col (out_col_17_5),
		.out_data (out_data_17_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_6;
	wire signed [DATA_WIDTH-1:0] out_col_17_6;
	wire signed [DATA_WIDTH-1:0] out_data_17_6;
	integer_mac_pe mac_pe_17_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_5),
		.in_col (out_col_16_6),
		.out_row (out_row_17_6),
		.out_col (out_col_17_6),
		.out_data (out_data_17_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_7;
	wire signed [DATA_WIDTH-1:0] out_col_17_7;
	wire signed [DATA_WIDTH-1:0] out_data_17_7;
	integer_mac_pe mac_pe_17_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_6),
		.in_col (out_col_16_7),
		.out_row (out_row_17_7),
		.out_col (out_col_17_7),
		.out_data (out_data_17_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_8;
	wire signed [DATA_WIDTH-1:0] out_col_17_8;
	wire signed [DATA_WIDTH-1:0] out_data_17_8;
	integer_mac_pe mac_pe_17_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_7),
		.in_col (out_col_16_8),
		.out_row (out_row_17_8),
		.out_col (out_col_17_8),
		.out_data (out_data_17_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_9;
	wire signed [DATA_WIDTH-1:0] out_col_17_9;
	wire signed [DATA_WIDTH-1:0] out_data_17_9;
	integer_mac_pe mac_pe_17_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_8),
		.in_col (out_col_16_9),
		.out_row (out_row_17_9),
		.out_col (out_col_17_9),
		.out_data (out_data_17_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_10;
	wire signed [DATA_WIDTH-1:0] out_col_17_10;
	wire signed [DATA_WIDTH-1:0] out_data_17_10;
	integer_mac_pe mac_pe_17_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_9),
		.in_col (out_col_16_10),
		.out_row (out_row_17_10),
		.out_col (out_col_17_10),
		.out_data (out_data_17_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_11;
	wire signed [DATA_WIDTH-1:0] out_col_17_11;
	wire signed [DATA_WIDTH-1:0] out_data_17_11;
	integer_mac_pe mac_pe_17_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_10),
		.in_col (out_col_16_11),
		.out_row (out_row_17_11),
		.out_col (out_col_17_11),
		.out_data (out_data_17_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_12;
	wire signed [DATA_WIDTH-1:0] out_col_17_12;
	wire signed [DATA_WIDTH-1:0] out_data_17_12;
	integer_mac_pe mac_pe_17_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_11),
		.in_col (out_col_16_12),
		.out_row (out_row_17_12),
		.out_col (out_col_17_12),
		.out_data (out_data_17_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_13;
	wire signed [DATA_WIDTH-1:0] out_col_17_13;
	wire signed [DATA_WIDTH-1:0] out_data_17_13;
	integer_mac_pe mac_pe_17_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_12),
		.in_col (out_col_16_13),
		.out_row (out_row_17_13),
		.out_col (out_col_17_13),
		.out_data (out_data_17_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_14;
	wire signed [DATA_WIDTH-1:0] out_col_17_14;
	wire signed [DATA_WIDTH-1:0] out_data_17_14;
	integer_mac_pe mac_pe_17_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_13),
		.in_col (out_col_16_14),
		.out_row (out_row_17_14),
		.out_col (out_col_17_14),
		.out_data (out_data_17_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_15;
	wire signed [DATA_WIDTH-1:0] out_col_17_15;
	wire signed [DATA_WIDTH-1:0] out_data_17_15;
	integer_mac_pe mac_pe_17_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_14),
		.in_col (out_col_16_15),
		.out_row (out_row_17_15),
		.out_col (out_col_17_15),
		.out_data (out_data_17_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_16;
	wire signed [DATA_WIDTH-1:0] out_col_17_16;
	wire signed [DATA_WIDTH-1:0] out_data_17_16;
	integer_mac_pe mac_pe_17_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_15),
		.in_col (out_col_16_16),
		.out_row (out_row_17_16),
		.out_col (out_col_17_16),
		.out_data (out_data_17_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_17;
	wire signed [DATA_WIDTH-1:0] out_col_17_17;
	wire signed [DATA_WIDTH-1:0] out_data_17_17;
	integer_mac_pe mac_pe_17_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_16),
		.in_col (out_col_16_17),
		.out_row (out_row_17_17),
		.out_col (out_col_17_17),
		.out_data (out_data_17_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_18;
	wire signed [DATA_WIDTH-1:0] out_col_17_18;
	wire signed [DATA_WIDTH-1:0] out_data_17_18;
	integer_mac_pe mac_pe_17_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_17),
		.in_col (out_col_16_18),
		.out_row (out_row_17_18),
		.out_col (out_col_17_18),
		.out_data (out_data_17_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_19;
	wire signed [DATA_WIDTH-1:0] out_col_17_19;
	wire signed [DATA_WIDTH-1:0] out_data_17_19;
	integer_mac_pe mac_pe_17_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_18),
		.in_col (out_col_16_19),
		.out_row (out_row_17_19),
		.out_col (out_col_17_19),
		.out_data (out_data_17_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_20;
	wire signed [DATA_WIDTH-1:0] out_col_17_20;
	wire signed [DATA_WIDTH-1:0] out_data_17_20;
	integer_mac_pe mac_pe_17_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_19),
		.in_col (out_col_16_20),
		.out_row (out_row_17_20),
		.out_col (out_col_17_20),
		.out_data (out_data_17_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_21;
	wire signed [DATA_WIDTH-1:0] out_col_17_21;
	wire signed [DATA_WIDTH-1:0] out_data_17_21;
	integer_mac_pe mac_pe_17_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_20),
		.in_col (out_col_16_21),
		.out_row (out_row_17_21),
		.out_col (out_col_17_21),
		.out_data (out_data_17_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_22;
	wire signed [DATA_WIDTH-1:0] out_col_17_22;
	wire signed [DATA_WIDTH-1:0] out_data_17_22;
	integer_mac_pe mac_pe_17_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_21),
		.in_col (out_col_16_22),
		.out_row (out_row_17_22),
		.out_col (out_col_17_22),
		.out_data (out_data_17_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_23;
	wire signed [DATA_WIDTH-1:0] out_col_17_23;
	wire signed [DATA_WIDTH-1:0] out_data_17_23;
	integer_mac_pe mac_pe_17_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_22),
		.in_col (out_col_16_23),
		.out_row (out_row_17_23),
		.out_col (out_col_17_23),
		.out_data (out_data_17_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_24;
	wire signed [DATA_WIDTH-1:0] out_col_17_24;
	wire signed [DATA_WIDTH-1:0] out_data_17_24;
	integer_mac_pe mac_pe_17_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_23),
		.in_col (out_col_16_24),
		.out_row (out_row_17_24),
		.out_col (out_col_17_24),
		.out_data (out_data_17_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_25;
	wire signed [DATA_WIDTH-1:0] out_col_17_25;
	wire signed [DATA_WIDTH-1:0] out_data_17_25;
	integer_mac_pe mac_pe_17_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_24),
		.in_col (out_col_16_25),
		.out_row (out_row_17_25),
		.out_col (out_col_17_25),
		.out_data (out_data_17_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_26;
	wire signed [DATA_WIDTH-1:0] out_col_17_26;
	wire signed [DATA_WIDTH-1:0] out_data_17_26;
	integer_mac_pe mac_pe_17_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_25),
		.in_col (out_col_16_26),
		.out_row (out_row_17_26),
		.out_col (out_col_17_26),
		.out_data (out_data_17_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_27;
	wire signed [DATA_WIDTH-1:0] out_col_17_27;
	wire signed [DATA_WIDTH-1:0] out_data_17_27;
	integer_mac_pe mac_pe_17_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_26),
		.in_col (out_col_16_27),
		.out_row (out_row_17_27),
		.out_col (out_col_17_27),
		.out_data (out_data_17_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_28;
	wire signed [DATA_WIDTH-1:0] out_col_17_28;
	wire signed [DATA_WIDTH-1:0] out_data_17_28;
	integer_mac_pe mac_pe_17_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_27),
		.in_col (out_col_16_28),
		.out_row (out_row_17_28),
		.out_col (out_col_17_28),
		.out_data (out_data_17_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_29;
	wire signed [DATA_WIDTH-1:0] out_col_17_29;
	wire signed [DATA_WIDTH-1:0] out_data_17_29;
	integer_mac_pe mac_pe_17_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_28),
		.in_col (out_col_16_29),
		.out_row (out_row_17_29),
		.out_col (out_col_17_29),
		.out_data (out_data_17_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_30;
	wire signed [DATA_WIDTH-1:0] out_col_17_30;
	wire signed [DATA_WIDTH-1:0] out_data_17_30;
	integer_mac_pe mac_pe_17_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_29),
		.in_col (out_col_16_30),
		.out_row (out_row_17_30),
		.out_col (out_col_17_30),
		.out_data (out_data_17_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_17_31;
	wire signed [DATA_WIDTH-1:0] out_col_17_31;
	wire signed [DATA_WIDTH-1:0] out_data_17_31;
	integer_mac_pe mac_pe_17_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_17_30),
		.in_col (out_col_16_31),
		.out_row (out_row_17_31),
		.out_col (out_col_17_31),
		.out_data (out_data_17_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_0;
	wire signed [DATA_WIDTH-1:0] out_col_18_0;
	wire signed [DATA_WIDTH-1:0] out_data_18_0;
	integer_mac_pe mac_pe_18_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_18_out),
		.in_col (out_col_17_0),
		.out_row (out_row_18_0),
		.out_col (out_col_18_0),
		.out_data (out_data_18_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_1;
	wire signed [DATA_WIDTH-1:0] out_col_18_1;
	wire signed [DATA_WIDTH-1:0] out_data_18_1;
	integer_mac_pe mac_pe_18_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_0),
		.in_col (out_col_17_1),
		.out_row (out_row_18_1),
		.out_col (out_col_18_1),
		.out_data (out_data_18_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_2;
	wire signed [DATA_WIDTH-1:0] out_col_18_2;
	wire signed [DATA_WIDTH-1:0] out_data_18_2;
	integer_mac_pe mac_pe_18_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_1),
		.in_col (out_col_17_2),
		.out_row (out_row_18_2),
		.out_col (out_col_18_2),
		.out_data (out_data_18_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_3;
	wire signed [DATA_WIDTH-1:0] out_col_18_3;
	wire signed [DATA_WIDTH-1:0] out_data_18_3;
	integer_mac_pe mac_pe_18_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_2),
		.in_col (out_col_17_3),
		.out_row (out_row_18_3),
		.out_col (out_col_18_3),
		.out_data (out_data_18_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_4;
	wire signed [DATA_WIDTH-1:0] out_col_18_4;
	wire signed [DATA_WIDTH-1:0] out_data_18_4;
	integer_mac_pe mac_pe_18_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_3),
		.in_col (out_col_17_4),
		.out_row (out_row_18_4),
		.out_col (out_col_18_4),
		.out_data (out_data_18_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_5;
	wire signed [DATA_WIDTH-1:0] out_col_18_5;
	wire signed [DATA_WIDTH-1:0] out_data_18_5;
	integer_mac_pe mac_pe_18_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_4),
		.in_col (out_col_17_5),
		.out_row (out_row_18_5),
		.out_col (out_col_18_5),
		.out_data (out_data_18_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_6;
	wire signed [DATA_WIDTH-1:0] out_col_18_6;
	wire signed [DATA_WIDTH-1:0] out_data_18_6;
	integer_mac_pe mac_pe_18_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_5),
		.in_col (out_col_17_6),
		.out_row (out_row_18_6),
		.out_col (out_col_18_6),
		.out_data (out_data_18_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_7;
	wire signed [DATA_WIDTH-1:0] out_col_18_7;
	wire signed [DATA_WIDTH-1:0] out_data_18_7;
	integer_mac_pe mac_pe_18_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_6),
		.in_col (out_col_17_7),
		.out_row (out_row_18_7),
		.out_col (out_col_18_7),
		.out_data (out_data_18_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_8;
	wire signed [DATA_WIDTH-1:0] out_col_18_8;
	wire signed [DATA_WIDTH-1:0] out_data_18_8;
	integer_mac_pe mac_pe_18_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_7),
		.in_col (out_col_17_8),
		.out_row (out_row_18_8),
		.out_col (out_col_18_8),
		.out_data (out_data_18_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_9;
	wire signed [DATA_WIDTH-1:0] out_col_18_9;
	wire signed [DATA_WIDTH-1:0] out_data_18_9;
	integer_mac_pe mac_pe_18_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_8),
		.in_col (out_col_17_9),
		.out_row (out_row_18_9),
		.out_col (out_col_18_9),
		.out_data (out_data_18_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_10;
	wire signed [DATA_WIDTH-1:0] out_col_18_10;
	wire signed [DATA_WIDTH-1:0] out_data_18_10;
	integer_mac_pe mac_pe_18_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_9),
		.in_col (out_col_17_10),
		.out_row (out_row_18_10),
		.out_col (out_col_18_10),
		.out_data (out_data_18_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_11;
	wire signed [DATA_WIDTH-1:0] out_col_18_11;
	wire signed [DATA_WIDTH-1:0] out_data_18_11;
	integer_mac_pe mac_pe_18_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_10),
		.in_col (out_col_17_11),
		.out_row (out_row_18_11),
		.out_col (out_col_18_11),
		.out_data (out_data_18_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_12;
	wire signed [DATA_WIDTH-1:0] out_col_18_12;
	wire signed [DATA_WIDTH-1:0] out_data_18_12;
	integer_mac_pe mac_pe_18_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_11),
		.in_col (out_col_17_12),
		.out_row (out_row_18_12),
		.out_col (out_col_18_12),
		.out_data (out_data_18_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_13;
	wire signed [DATA_WIDTH-1:0] out_col_18_13;
	wire signed [DATA_WIDTH-1:0] out_data_18_13;
	integer_mac_pe mac_pe_18_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_12),
		.in_col (out_col_17_13),
		.out_row (out_row_18_13),
		.out_col (out_col_18_13),
		.out_data (out_data_18_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_14;
	wire signed [DATA_WIDTH-1:0] out_col_18_14;
	wire signed [DATA_WIDTH-1:0] out_data_18_14;
	integer_mac_pe mac_pe_18_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_13),
		.in_col (out_col_17_14),
		.out_row (out_row_18_14),
		.out_col (out_col_18_14),
		.out_data (out_data_18_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_15;
	wire signed [DATA_WIDTH-1:0] out_col_18_15;
	wire signed [DATA_WIDTH-1:0] out_data_18_15;
	integer_mac_pe mac_pe_18_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_14),
		.in_col (out_col_17_15),
		.out_row (out_row_18_15),
		.out_col (out_col_18_15),
		.out_data (out_data_18_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_16;
	wire signed [DATA_WIDTH-1:0] out_col_18_16;
	wire signed [DATA_WIDTH-1:0] out_data_18_16;
	integer_mac_pe mac_pe_18_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_15),
		.in_col (out_col_17_16),
		.out_row (out_row_18_16),
		.out_col (out_col_18_16),
		.out_data (out_data_18_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_17;
	wire signed [DATA_WIDTH-1:0] out_col_18_17;
	wire signed [DATA_WIDTH-1:0] out_data_18_17;
	integer_mac_pe mac_pe_18_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_16),
		.in_col (out_col_17_17),
		.out_row (out_row_18_17),
		.out_col (out_col_18_17),
		.out_data (out_data_18_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_18;
	wire signed [DATA_WIDTH-1:0] out_col_18_18;
	wire signed [DATA_WIDTH-1:0] out_data_18_18;
	integer_mac_pe mac_pe_18_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_17),
		.in_col (out_col_17_18),
		.out_row (out_row_18_18),
		.out_col (out_col_18_18),
		.out_data (out_data_18_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_19;
	wire signed [DATA_WIDTH-1:0] out_col_18_19;
	wire signed [DATA_WIDTH-1:0] out_data_18_19;
	integer_mac_pe mac_pe_18_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_18),
		.in_col (out_col_17_19),
		.out_row (out_row_18_19),
		.out_col (out_col_18_19),
		.out_data (out_data_18_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_20;
	wire signed [DATA_WIDTH-1:0] out_col_18_20;
	wire signed [DATA_WIDTH-1:0] out_data_18_20;
	integer_mac_pe mac_pe_18_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_19),
		.in_col (out_col_17_20),
		.out_row (out_row_18_20),
		.out_col (out_col_18_20),
		.out_data (out_data_18_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_21;
	wire signed [DATA_WIDTH-1:0] out_col_18_21;
	wire signed [DATA_WIDTH-1:0] out_data_18_21;
	integer_mac_pe mac_pe_18_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_20),
		.in_col (out_col_17_21),
		.out_row (out_row_18_21),
		.out_col (out_col_18_21),
		.out_data (out_data_18_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_22;
	wire signed [DATA_WIDTH-1:0] out_col_18_22;
	wire signed [DATA_WIDTH-1:0] out_data_18_22;
	integer_mac_pe mac_pe_18_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_21),
		.in_col (out_col_17_22),
		.out_row (out_row_18_22),
		.out_col (out_col_18_22),
		.out_data (out_data_18_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_23;
	wire signed [DATA_WIDTH-1:0] out_col_18_23;
	wire signed [DATA_WIDTH-1:0] out_data_18_23;
	integer_mac_pe mac_pe_18_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_22),
		.in_col (out_col_17_23),
		.out_row (out_row_18_23),
		.out_col (out_col_18_23),
		.out_data (out_data_18_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_24;
	wire signed [DATA_WIDTH-1:0] out_col_18_24;
	wire signed [DATA_WIDTH-1:0] out_data_18_24;
	integer_mac_pe mac_pe_18_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_23),
		.in_col (out_col_17_24),
		.out_row (out_row_18_24),
		.out_col (out_col_18_24),
		.out_data (out_data_18_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_25;
	wire signed [DATA_WIDTH-1:0] out_col_18_25;
	wire signed [DATA_WIDTH-1:0] out_data_18_25;
	integer_mac_pe mac_pe_18_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_24),
		.in_col (out_col_17_25),
		.out_row (out_row_18_25),
		.out_col (out_col_18_25),
		.out_data (out_data_18_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_26;
	wire signed [DATA_WIDTH-1:0] out_col_18_26;
	wire signed [DATA_WIDTH-1:0] out_data_18_26;
	integer_mac_pe mac_pe_18_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_25),
		.in_col (out_col_17_26),
		.out_row (out_row_18_26),
		.out_col (out_col_18_26),
		.out_data (out_data_18_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_27;
	wire signed [DATA_WIDTH-1:0] out_col_18_27;
	wire signed [DATA_WIDTH-1:0] out_data_18_27;
	integer_mac_pe mac_pe_18_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_26),
		.in_col (out_col_17_27),
		.out_row (out_row_18_27),
		.out_col (out_col_18_27),
		.out_data (out_data_18_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_28;
	wire signed [DATA_WIDTH-1:0] out_col_18_28;
	wire signed [DATA_WIDTH-1:0] out_data_18_28;
	integer_mac_pe mac_pe_18_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_27),
		.in_col (out_col_17_28),
		.out_row (out_row_18_28),
		.out_col (out_col_18_28),
		.out_data (out_data_18_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_29;
	wire signed [DATA_WIDTH-1:0] out_col_18_29;
	wire signed [DATA_WIDTH-1:0] out_data_18_29;
	integer_mac_pe mac_pe_18_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_28),
		.in_col (out_col_17_29),
		.out_row (out_row_18_29),
		.out_col (out_col_18_29),
		.out_data (out_data_18_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_30;
	wire signed [DATA_WIDTH-1:0] out_col_18_30;
	wire signed [DATA_WIDTH-1:0] out_data_18_30;
	integer_mac_pe mac_pe_18_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_29),
		.in_col (out_col_17_30),
		.out_row (out_row_18_30),
		.out_col (out_col_18_30),
		.out_data (out_data_18_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_18_31;
	wire signed [DATA_WIDTH-1:0] out_col_18_31;
	wire signed [DATA_WIDTH-1:0] out_data_18_31;
	integer_mac_pe mac_pe_18_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_18_30),
		.in_col (out_col_17_31),
		.out_row (out_row_18_31),
		.out_col (out_col_18_31),
		.out_data (out_data_18_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_0;
	wire signed [DATA_WIDTH-1:0] out_col_19_0;
	wire signed [DATA_WIDTH-1:0] out_data_19_0;
	integer_mac_pe mac_pe_19_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_19_out),
		.in_col (out_col_18_0),
		.out_row (out_row_19_0),
		.out_col (out_col_19_0),
		.out_data (out_data_19_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_1;
	wire signed [DATA_WIDTH-1:0] out_col_19_1;
	wire signed [DATA_WIDTH-1:0] out_data_19_1;
	integer_mac_pe mac_pe_19_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_0),
		.in_col (out_col_18_1),
		.out_row (out_row_19_1),
		.out_col (out_col_19_1),
		.out_data (out_data_19_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_2;
	wire signed [DATA_WIDTH-1:0] out_col_19_2;
	wire signed [DATA_WIDTH-1:0] out_data_19_2;
	integer_mac_pe mac_pe_19_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_1),
		.in_col (out_col_18_2),
		.out_row (out_row_19_2),
		.out_col (out_col_19_2),
		.out_data (out_data_19_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_3;
	wire signed [DATA_WIDTH-1:0] out_col_19_3;
	wire signed [DATA_WIDTH-1:0] out_data_19_3;
	integer_mac_pe mac_pe_19_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_2),
		.in_col (out_col_18_3),
		.out_row (out_row_19_3),
		.out_col (out_col_19_3),
		.out_data (out_data_19_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_4;
	wire signed [DATA_WIDTH-1:0] out_col_19_4;
	wire signed [DATA_WIDTH-1:0] out_data_19_4;
	integer_mac_pe mac_pe_19_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_3),
		.in_col (out_col_18_4),
		.out_row (out_row_19_4),
		.out_col (out_col_19_4),
		.out_data (out_data_19_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_5;
	wire signed [DATA_WIDTH-1:0] out_col_19_5;
	wire signed [DATA_WIDTH-1:0] out_data_19_5;
	integer_mac_pe mac_pe_19_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_4),
		.in_col (out_col_18_5),
		.out_row (out_row_19_5),
		.out_col (out_col_19_5),
		.out_data (out_data_19_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_6;
	wire signed [DATA_WIDTH-1:0] out_col_19_6;
	wire signed [DATA_WIDTH-1:0] out_data_19_6;
	integer_mac_pe mac_pe_19_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_5),
		.in_col (out_col_18_6),
		.out_row (out_row_19_6),
		.out_col (out_col_19_6),
		.out_data (out_data_19_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_7;
	wire signed [DATA_WIDTH-1:0] out_col_19_7;
	wire signed [DATA_WIDTH-1:0] out_data_19_7;
	integer_mac_pe mac_pe_19_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_6),
		.in_col (out_col_18_7),
		.out_row (out_row_19_7),
		.out_col (out_col_19_7),
		.out_data (out_data_19_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_8;
	wire signed [DATA_WIDTH-1:0] out_col_19_8;
	wire signed [DATA_WIDTH-1:0] out_data_19_8;
	integer_mac_pe mac_pe_19_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_7),
		.in_col (out_col_18_8),
		.out_row (out_row_19_8),
		.out_col (out_col_19_8),
		.out_data (out_data_19_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_9;
	wire signed [DATA_WIDTH-1:0] out_col_19_9;
	wire signed [DATA_WIDTH-1:0] out_data_19_9;
	integer_mac_pe mac_pe_19_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_8),
		.in_col (out_col_18_9),
		.out_row (out_row_19_9),
		.out_col (out_col_19_9),
		.out_data (out_data_19_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_10;
	wire signed [DATA_WIDTH-1:0] out_col_19_10;
	wire signed [DATA_WIDTH-1:0] out_data_19_10;
	integer_mac_pe mac_pe_19_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_9),
		.in_col (out_col_18_10),
		.out_row (out_row_19_10),
		.out_col (out_col_19_10),
		.out_data (out_data_19_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_11;
	wire signed [DATA_WIDTH-1:0] out_col_19_11;
	wire signed [DATA_WIDTH-1:0] out_data_19_11;
	integer_mac_pe mac_pe_19_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_10),
		.in_col (out_col_18_11),
		.out_row (out_row_19_11),
		.out_col (out_col_19_11),
		.out_data (out_data_19_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_12;
	wire signed [DATA_WIDTH-1:0] out_col_19_12;
	wire signed [DATA_WIDTH-1:0] out_data_19_12;
	integer_mac_pe mac_pe_19_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_11),
		.in_col (out_col_18_12),
		.out_row (out_row_19_12),
		.out_col (out_col_19_12),
		.out_data (out_data_19_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_13;
	wire signed [DATA_WIDTH-1:0] out_col_19_13;
	wire signed [DATA_WIDTH-1:0] out_data_19_13;
	integer_mac_pe mac_pe_19_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_12),
		.in_col (out_col_18_13),
		.out_row (out_row_19_13),
		.out_col (out_col_19_13),
		.out_data (out_data_19_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_14;
	wire signed [DATA_WIDTH-1:0] out_col_19_14;
	wire signed [DATA_WIDTH-1:0] out_data_19_14;
	integer_mac_pe mac_pe_19_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_13),
		.in_col (out_col_18_14),
		.out_row (out_row_19_14),
		.out_col (out_col_19_14),
		.out_data (out_data_19_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_15;
	wire signed [DATA_WIDTH-1:0] out_col_19_15;
	wire signed [DATA_WIDTH-1:0] out_data_19_15;
	integer_mac_pe mac_pe_19_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_14),
		.in_col (out_col_18_15),
		.out_row (out_row_19_15),
		.out_col (out_col_19_15),
		.out_data (out_data_19_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_16;
	wire signed [DATA_WIDTH-1:0] out_col_19_16;
	wire signed [DATA_WIDTH-1:0] out_data_19_16;
	integer_mac_pe mac_pe_19_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_15),
		.in_col (out_col_18_16),
		.out_row (out_row_19_16),
		.out_col (out_col_19_16),
		.out_data (out_data_19_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_17;
	wire signed [DATA_WIDTH-1:0] out_col_19_17;
	wire signed [DATA_WIDTH-1:0] out_data_19_17;
	integer_mac_pe mac_pe_19_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_16),
		.in_col (out_col_18_17),
		.out_row (out_row_19_17),
		.out_col (out_col_19_17),
		.out_data (out_data_19_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_18;
	wire signed [DATA_WIDTH-1:0] out_col_19_18;
	wire signed [DATA_WIDTH-1:0] out_data_19_18;
	integer_mac_pe mac_pe_19_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_17),
		.in_col (out_col_18_18),
		.out_row (out_row_19_18),
		.out_col (out_col_19_18),
		.out_data (out_data_19_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_19;
	wire signed [DATA_WIDTH-1:0] out_col_19_19;
	wire signed [DATA_WIDTH-1:0] out_data_19_19;
	integer_mac_pe mac_pe_19_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_18),
		.in_col (out_col_18_19),
		.out_row (out_row_19_19),
		.out_col (out_col_19_19),
		.out_data (out_data_19_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_20;
	wire signed [DATA_WIDTH-1:0] out_col_19_20;
	wire signed [DATA_WIDTH-1:0] out_data_19_20;
	integer_mac_pe mac_pe_19_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_19),
		.in_col (out_col_18_20),
		.out_row (out_row_19_20),
		.out_col (out_col_19_20),
		.out_data (out_data_19_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_21;
	wire signed [DATA_WIDTH-1:0] out_col_19_21;
	wire signed [DATA_WIDTH-1:0] out_data_19_21;
	integer_mac_pe mac_pe_19_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_20),
		.in_col (out_col_18_21),
		.out_row (out_row_19_21),
		.out_col (out_col_19_21),
		.out_data (out_data_19_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_22;
	wire signed [DATA_WIDTH-1:0] out_col_19_22;
	wire signed [DATA_WIDTH-1:0] out_data_19_22;
	integer_mac_pe mac_pe_19_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_21),
		.in_col (out_col_18_22),
		.out_row (out_row_19_22),
		.out_col (out_col_19_22),
		.out_data (out_data_19_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_23;
	wire signed [DATA_WIDTH-1:0] out_col_19_23;
	wire signed [DATA_WIDTH-1:0] out_data_19_23;
	integer_mac_pe mac_pe_19_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_22),
		.in_col (out_col_18_23),
		.out_row (out_row_19_23),
		.out_col (out_col_19_23),
		.out_data (out_data_19_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_24;
	wire signed [DATA_WIDTH-1:0] out_col_19_24;
	wire signed [DATA_WIDTH-1:0] out_data_19_24;
	integer_mac_pe mac_pe_19_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_23),
		.in_col (out_col_18_24),
		.out_row (out_row_19_24),
		.out_col (out_col_19_24),
		.out_data (out_data_19_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_25;
	wire signed [DATA_WIDTH-1:0] out_col_19_25;
	wire signed [DATA_WIDTH-1:0] out_data_19_25;
	integer_mac_pe mac_pe_19_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_24),
		.in_col (out_col_18_25),
		.out_row (out_row_19_25),
		.out_col (out_col_19_25),
		.out_data (out_data_19_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_26;
	wire signed [DATA_WIDTH-1:0] out_col_19_26;
	wire signed [DATA_WIDTH-1:0] out_data_19_26;
	integer_mac_pe mac_pe_19_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_25),
		.in_col (out_col_18_26),
		.out_row (out_row_19_26),
		.out_col (out_col_19_26),
		.out_data (out_data_19_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_27;
	wire signed [DATA_WIDTH-1:0] out_col_19_27;
	wire signed [DATA_WIDTH-1:0] out_data_19_27;
	integer_mac_pe mac_pe_19_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_26),
		.in_col (out_col_18_27),
		.out_row (out_row_19_27),
		.out_col (out_col_19_27),
		.out_data (out_data_19_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_28;
	wire signed [DATA_WIDTH-1:0] out_col_19_28;
	wire signed [DATA_WIDTH-1:0] out_data_19_28;
	integer_mac_pe mac_pe_19_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_27),
		.in_col (out_col_18_28),
		.out_row (out_row_19_28),
		.out_col (out_col_19_28),
		.out_data (out_data_19_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_29;
	wire signed [DATA_WIDTH-1:0] out_col_19_29;
	wire signed [DATA_WIDTH-1:0] out_data_19_29;
	integer_mac_pe mac_pe_19_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_28),
		.in_col (out_col_18_29),
		.out_row (out_row_19_29),
		.out_col (out_col_19_29),
		.out_data (out_data_19_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_30;
	wire signed [DATA_WIDTH-1:0] out_col_19_30;
	wire signed [DATA_WIDTH-1:0] out_data_19_30;
	integer_mac_pe mac_pe_19_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_29),
		.in_col (out_col_18_30),
		.out_row (out_row_19_30),
		.out_col (out_col_19_30),
		.out_data (out_data_19_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_19_31;
	wire signed [DATA_WIDTH-1:0] out_col_19_31;
	wire signed [DATA_WIDTH-1:0] out_data_19_31;
	integer_mac_pe mac_pe_19_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_19_30),
		.in_col (out_col_18_31),
		.out_row (out_row_19_31),
		.out_col (out_col_19_31),
		.out_data (out_data_19_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_0;
	wire signed [DATA_WIDTH-1:0] out_col_20_0;
	wire signed [DATA_WIDTH-1:0] out_data_20_0;
	integer_mac_pe mac_pe_20_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_20_out),
		.in_col (out_col_19_0),
		.out_row (out_row_20_0),
		.out_col (out_col_20_0),
		.out_data (out_data_20_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_1;
	wire signed [DATA_WIDTH-1:0] out_col_20_1;
	wire signed [DATA_WIDTH-1:0] out_data_20_1;
	integer_mac_pe mac_pe_20_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_0),
		.in_col (out_col_19_1),
		.out_row (out_row_20_1),
		.out_col (out_col_20_1),
		.out_data (out_data_20_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_2;
	wire signed [DATA_WIDTH-1:0] out_col_20_2;
	wire signed [DATA_WIDTH-1:0] out_data_20_2;
	integer_mac_pe mac_pe_20_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_1),
		.in_col (out_col_19_2),
		.out_row (out_row_20_2),
		.out_col (out_col_20_2),
		.out_data (out_data_20_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_3;
	wire signed [DATA_WIDTH-1:0] out_col_20_3;
	wire signed [DATA_WIDTH-1:0] out_data_20_3;
	integer_mac_pe mac_pe_20_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_2),
		.in_col (out_col_19_3),
		.out_row (out_row_20_3),
		.out_col (out_col_20_3),
		.out_data (out_data_20_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_4;
	wire signed [DATA_WIDTH-1:0] out_col_20_4;
	wire signed [DATA_WIDTH-1:0] out_data_20_4;
	integer_mac_pe mac_pe_20_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_3),
		.in_col (out_col_19_4),
		.out_row (out_row_20_4),
		.out_col (out_col_20_4),
		.out_data (out_data_20_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_5;
	wire signed [DATA_WIDTH-1:0] out_col_20_5;
	wire signed [DATA_WIDTH-1:0] out_data_20_5;
	integer_mac_pe mac_pe_20_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_4),
		.in_col (out_col_19_5),
		.out_row (out_row_20_5),
		.out_col (out_col_20_5),
		.out_data (out_data_20_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_6;
	wire signed [DATA_WIDTH-1:0] out_col_20_6;
	wire signed [DATA_WIDTH-1:0] out_data_20_6;
	integer_mac_pe mac_pe_20_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_5),
		.in_col (out_col_19_6),
		.out_row (out_row_20_6),
		.out_col (out_col_20_6),
		.out_data (out_data_20_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_7;
	wire signed [DATA_WIDTH-1:0] out_col_20_7;
	wire signed [DATA_WIDTH-1:0] out_data_20_7;
	integer_mac_pe mac_pe_20_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_6),
		.in_col (out_col_19_7),
		.out_row (out_row_20_7),
		.out_col (out_col_20_7),
		.out_data (out_data_20_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_8;
	wire signed [DATA_WIDTH-1:0] out_col_20_8;
	wire signed [DATA_WIDTH-1:0] out_data_20_8;
	integer_mac_pe mac_pe_20_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_7),
		.in_col (out_col_19_8),
		.out_row (out_row_20_8),
		.out_col (out_col_20_8),
		.out_data (out_data_20_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_9;
	wire signed [DATA_WIDTH-1:0] out_col_20_9;
	wire signed [DATA_WIDTH-1:0] out_data_20_9;
	integer_mac_pe mac_pe_20_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_8),
		.in_col (out_col_19_9),
		.out_row (out_row_20_9),
		.out_col (out_col_20_9),
		.out_data (out_data_20_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_10;
	wire signed [DATA_WIDTH-1:0] out_col_20_10;
	wire signed [DATA_WIDTH-1:0] out_data_20_10;
	integer_mac_pe mac_pe_20_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_9),
		.in_col (out_col_19_10),
		.out_row (out_row_20_10),
		.out_col (out_col_20_10),
		.out_data (out_data_20_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_11;
	wire signed [DATA_WIDTH-1:0] out_col_20_11;
	wire signed [DATA_WIDTH-1:0] out_data_20_11;
	integer_mac_pe mac_pe_20_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_10),
		.in_col (out_col_19_11),
		.out_row (out_row_20_11),
		.out_col (out_col_20_11),
		.out_data (out_data_20_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_12;
	wire signed [DATA_WIDTH-1:0] out_col_20_12;
	wire signed [DATA_WIDTH-1:0] out_data_20_12;
	integer_mac_pe mac_pe_20_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_11),
		.in_col (out_col_19_12),
		.out_row (out_row_20_12),
		.out_col (out_col_20_12),
		.out_data (out_data_20_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_13;
	wire signed [DATA_WIDTH-1:0] out_col_20_13;
	wire signed [DATA_WIDTH-1:0] out_data_20_13;
	integer_mac_pe mac_pe_20_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_12),
		.in_col (out_col_19_13),
		.out_row (out_row_20_13),
		.out_col (out_col_20_13),
		.out_data (out_data_20_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_14;
	wire signed [DATA_WIDTH-1:0] out_col_20_14;
	wire signed [DATA_WIDTH-1:0] out_data_20_14;
	integer_mac_pe mac_pe_20_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_13),
		.in_col (out_col_19_14),
		.out_row (out_row_20_14),
		.out_col (out_col_20_14),
		.out_data (out_data_20_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_15;
	wire signed [DATA_WIDTH-1:0] out_col_20_15;
	wire signed [DATA_WIDTH-1:0] out_data_20_15;
	integer_mac_pe mac_pe_20_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_14),
		.in_col (out_col_19_15),
		.out_row (out_row_20_15),
		.out_col (out_col_20_15),
		.out_data (out_data_20_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_16;
	wire signed [DATA_WIDTH-1:0] out_col_20_16;
	wire signed [DATA_WIDTH-1:0] out_data_20_16;
	integer_mac_pe mac_pe_20_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_15),
		.in_col (out_col_19_16),
		.out_row (out_row_20_16),
		.out_col (out_col_20_16),
		.out_data (out_data_20_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_17;
	wire signed [DATA_WIDTH-1:0] out_col_20_17;
	wire signed [DATA_WIDTH-1:0] out_data_20_17;
	integer_mac_pe mac_pe_20_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_16),
		.in_col (out_col_19_17),
		.out_row (out_row_20_17),
		.out_col (out_col_20_17),
		.out_data (out_data_20_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_18;
	wire signed [DATA_WIDTH-1:0] out_col_20_18;
	wire signed [DATA_WIDTH-1:0] out_data_20_18;
	integer_mac_pe mac_pe_20_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_17),
		.in_col (out_col_19_18),
		.out_row (out_row_20_18),
		.out_col (out_col_20_18),
		.out_data (out_data_20_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_19;
	wire signed [DATA_WIDTH-1:0] out_col_20_19;
	wire signed [DATA_WIDTH-1:0] out_data_20_19;
	integer_mac_pe mac_pe_20_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_18),
		.in_col (out_col_19_19),
		.out_row (out_row_20_19),
		.out_col (out_col_20_19),
		.out_data (out_data_20_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_20;
	wire signed [DATA_WIDTH-1:0] out_col_20_20;
	wire signed [DATA_WIDTH-1:0] out_data_20_20;
	integer_mac_pe mac_pe_20_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_19),
		.in_col (out_col_19_20),
		.out_row (out_row_20_20),
		.out_col (out_col_20_20),
		.out_data (out_data_20_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_21;
	wire signed [DATA_WIDTH-1:0] out_col_20_21;
	wire signed [DATA_WIDTH-1:0] out_data_20_21;
	integer_mac_pe mac_pe_20_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_20),
		.in_col (out_col_19_21),
		.out_row (out_row_20_21),
		.out_col (out_col_20_21),
		.out_data (out_data_20_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_22;
	wire signed [DATA_WIDTH-1:0] out_col_20_22;
	wire signed [DATA_WIDTH-1:0] out_data_20_22;
	integer_mac_pe mac_pe_20_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_21),
		.in_col (out_col_19_22),
		.out_row (out_row_20_22),
		.out_col (out_col_20_22),
		.out_data (out_data_20_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_23;
	wire signed [DATA_WIDTH-1:0] out_col_20_23;
	wire signed [DATA_WIDTH-1:0] out_data_20_23;
	integer_mac_pe mac_pe_20_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_22),
		.in_col (out_col_19_23),
		.out_row (out_row_20_23),
		.out_col (out_col_20_23),
		.out_data (out_data_20_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_24;
	wire signed [DATA_WIDTH-1:0] out_col_20_24;
	wire signed [DATA_WIDTH-1:0] out_data_20_24;
	integer_mac_pe mac_pe_20_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_23),
		.in_col (out_col_19_24),
		.out_row (out_row_20_24),
		.out_col (out_col_20_24),
		.out_data (out_data_20_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_25;
	wire signed [DATA_WIDTH-1:0] out_col_20_25;
	wire signed [DATA_WIDTH-1:0] out_data_20_25;
	integer_mac_pe mac_pe_20_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_24),
		.in_col (out_col_19_25),
		.out_row (out_row_20_25),
		.out_col (out_col_20_25),
		.out_data (out_data_20_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_26;
	wire signed [DATA_WIDTH-1:0] out_col_20_26;
	wire signed [DATA_WIDTH-1:0] out_data_20_26;
	integer_mac_pe mac_pe_20_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_25),
		.in_col (out_col_19_26),
		.out_row (out_row_20_26),
		.out_col (out_col_20_26),
		.out_data (out_data_20_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_27;
	wire signed [DATA_WIDTH-1:0] out_col_20_27;
	wire signed [DATA_WIDTH-1:0] out_data_20_27;
	integer_mac_pe mac_pe_20_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_26),
		.in_col (out_col_19_27),
		.out_row (out_row_20_27),
		.out_col (out_col_20_27),
		.out_data (out_data_20_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_28;
	wire signed [DATA_WIDTH-1:0] out_col_20_28;
	wire signed [DATA_WIDTH-1:0] out_data_20_28;
	integer_mac_pe mac_pe_20_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_27),
		.in_col (out_col_19_28),
		.out_row (out_row_20_28),
		.out_col (out_col_20_28),
		.out_data (out_data_20_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_29;
	wire signed [DATA_WIDTH-1:0] out_col_20_29;
	wire signed [DATA_WIDTH-1:0] out_data_20_29;
	integer_mac_pe mac_pe_20_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_28),
		.in_col (out_col_19_29),
		.out_row (out_row_20_29),
		.out_col (out_col_20_29),
		.out_data (out_data_20_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_30;
	wire signed [DATA_WIDTH-1:0] out_col_20_30;
	wire signed [DATA_WIDTH-1:0] out_data_20_30;
	integer_mac_pe mac_pe_20_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_29),
		.in_col (out_col_19_30),
		.out_row (out_row_20_30),
		.out_col (out_col_20_30),
		.out_data (out_data_20_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_20_31;
	wire signed [DATA_WIDTH-1:0] out_col_20_31;
	wire signed [DATA_WIDTH-1:0] out_data_20_31;
	integer_mac_pe mac_pe_20_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_20_30),
		.in_col (out_col_19_31),
		.out_row (out_row_20_31),
		.out_col (out_col_20_31),
		.out_data (out_data_20_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_0;
	wire signed [DATA_WIDTH-1:0] out_col_21_0;
	wire signed [DATA_WIDTH-1:0] out_data_21_0;
	integer_mac_pe mac_pe_21_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_21_out),
		.in_col (out_col_20_0),
		.out_row (out_row_21_0),
		.out_col (out_col_21_0),
		.out_data (out_data_21_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_1;
	wire signed [DATA_WIDTH-1:0] out_col_21_1;
	wire signed [DATA_WIDTH-1:0] out_data_21_1;
	integer_mac_pe mac_pe_21_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_0),
		.in_col (out_col_20_1),
		.out_row (out_row_21_1),
		.out_col (out_col_21_1),
		.out_data (out_data_21_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_2;
	wire signed [DATA_WIDTH-1:0] out_col_21_2;
	wire signed [DATA_WIDTH-1:0] out_data_21_2;
	integer_mac_pe mac_pe_21_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_1),
		.in_col (out_col_20_2),
		.out_row (out_row_21_2),
		.out_col (out_col_21_2),
		.out_data (out_data_21_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_3;
	wire signed [DATA_WIDTH-1:0] out_col_21_3;
	wire signed [DATA_WIDTH-1:0] out_data_21_3;
	integer_mac_pe mac_pe_21_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_2),
		.in_col (out_col_20_3),
		.out_row (out_row_21_3),
		.out_col (out_col_21_3),
		.out_data (out_data_21_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_4;
	wire signed [DATA_WIDTH-1:0] out_col_21_4;
	wire signed [DATA_WIDTH-1:0] out_data_21_4;
	integer_mac_pe mac_pe_21_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_3),
		.in_col (out_col_20_4),
		.out_row (out_row_21_4),
		.out_col (out_col_21_4),
		.out_data (out_data_21_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_5;
	wire signed [DATA_WIDTH-1:0] out_col_21_5;
	wire signed [DATA_WIDTH-1:0] out_data_21_5;
	integer_mac_pe mac_pe_21_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_4),
		.in_col (out_col_20_5),
		.out_row (out_row_21_5),
		.out_col (out_col_21_5),
		.out_data (out_data_21_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_6;
	wire signed [DATA_WIDTH-1:0] out_col_21_6;
	wire signed [DATA_WIDTH-1:0] out_data_21_6;
	integer_mac_pe mac_pe_21_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_5),
		.in_col (out_col_20_6),
		.out_row (out_row_21_6),
		.out_col (out_col_21_6),
		.out_data (out_data_21_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_7;
	wire signed [DATA_WIDTH-1:0] out_col_21_7;
	wire signed [DATA_WIDTH-1:0] out_data_21_7;
	integer_mac_pe mac_pe_21_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_6),
		.in_col (out_col_20_7),
		.out_row (out_row_21_7),
		.out_col (out_col_21_7),
		.out_data (out_data_21_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_8;
	wire signed [DATA_WIDTH-1:0] out_col_21_8;
	wire signed [DATA_WIDTH-1:0] out_data_21_8;
	integer_mac_pe mac_pe_21_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_7),
		.in_col (out_col_20_8),
		.out_row (out_row_21_8),
		.out_col (out_col_21_8),
		.out_data (out_data_21_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_9;
	wire signed [DATA_WIDTH-1:0] out_col_21_9;
	wire signed [DATA_WIDTH-1:0] out_data_21_9;
	integer_mac_pe mac_pe_21_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_8),
		.in_col (out_col_20_9),
		.out_row (out_row_21_9),
		.out_col (out_col_21_9),
		.out_data (out_data_21_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_10;
	wire signed [DATA_WIDTH-1:0] out_col_21_10;
	wire signed [DATA_WIDTH-1:0] out_data_21_10;
	integer_mac_pe mac_pe_21_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_9),
		.in_col (out_col_20_10),
		.out_row (out_row_21_10),
		.out_col (out_col_21_10),
		.out_data (out_data_21_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_11;
	wire signed [DATA_WIDTH-1:0] out_col_21_11;
	wire signed [DATA_WIDTH-1:0] out_data_21_11;
	integer_mac_pe mac_pe_21_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_10),
		.in_col (out_col_20_11),
		.out_row (out_row_21_11),
		.out_col (out_col_21_11),
		.out_data (out_data_21_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_12;
	wire signed [DATA_WIDTH-1:0] out_col_21_12;
	wire signed [DATA_WIDTH-1:0] out_data_21_12;
	integer_mac_pe mac_pe_21_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_11),
		.in_col (out_col_20_12),
		.out_row (out_row_21_12),
		.out_col (out_col_21_12),
		.out_data (out_data_21_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_13;
	wire signed [DATA_WIDTH-1:0] out_col_21_13;
	wire signed [DATA_WIDTH-1:0] out_data_21_13;
	integer_mac_pe mac_pe_21_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_12),
		.in_col (out_col_20_13),
		.out_row (out_row_21_13),
		.out_col (out_col_21_13),
		.out_data (out_data_21_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_14;
	wire signed [DATA_WIDTH-1:0] out_col_21_14;
	wire signed [DATA_WIDTH-1:0] out_data_21_14;
	integer_mac_pe mac_pe_21_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_13),
		.in_col (out_col_20_14),
		.out_row (out_row_21_14),
		.out_col (out_col_21_14),
		.out_data (out_data_21_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_15;
	wire signed [DATA_WIDTH-1:0] out_col_21_15;
	wire signed [DATA_WIDTH-1:0] out_data_21_15;
	integer_mac_pe mac_pe_21_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_14),
		.in_col (out_col_20_15),
		.out_row (out_row_21_15),
		.out_col (out_col_21_15),
		.out_data (out_data_21_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_16;
	wire signed [DATA_WIDTH-1:0] out_col_21_16;
	wire signed [DATA_WIDTH-1:0] out_data_21_16;
	integer_mac_pe mac_pe_21_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_15),
		.in_col (out_col_20_16),
		.out_row (out_row_21_16),
		.out_col (out_col_21_16),
		.out_data (out_data_21_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_17;
	wire signed [DATA_WIDTH-1:0] out_col_21_17;
	wire signed [DATA_WIDTH-1:0] out_data_21_17;
	integer_mac_pe mac_pe_21_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_16),
		.in_col (out_col_20_17),
		.out_row (out_row_21_17),
		.out_col (out_col_21_17),
		.out_data (out_data_21_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_18;
	wire signed [DATA_WIDTH-1:0] out_col_21_18;
	wire signed [DATA_WIDTH-1:0] out_data_21_18;
	integer_mac_pe mac_pe_21_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_17),
		.in_col (out_col_20_18),
		.out_row (out_row_21_18),
		.out_col (out_col_21_18),
		.out_data (out_data_21_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_19;
	wire signed [DATA_WIDTH-1:0] out_col_21_19;
	wire signed [DATA_WIDTH-1:0] out_data_21_19;
	integer_mac_pe mac_pe_21_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_18),
		.in_col (out_col_20_19),
		.out_row (out_row_21_19),
		.out_col (out_col_21_19),
		.out_data (out_data_21_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_20;
	wire signed [DATA_WIDTH-1:0] out_col_21_20;
	wire signed [DATA_WIDTH-1:0] out_data_21_20;
	integer_mac_pe mac_pe_21_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_19),
		.in_col (out_col_20_20),
		.out_row (out_row_21_20),
		.out_col (out_col_21_20),
		.out_data (out_data_21_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_21;
	wire signed [DATA_WIDTH-1:0] out_col_21_21;
	wire signed [DATA_WIDTH-1:0] out_data_21_21;
	integer_mac_pe mac_pe_21_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_20),
		.in_col (out_col_20_21),
		.out_row (out_row_21_21),
		.out_col (out_col_21_21),
		.out_data (out_data_21_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_22;
	wire signed [DATA_WIDTH-1:0] out_col_21_22;
	wire signed [DATA_WIDTH-1:0] out_data_21_22;
	integer_mac_pe mac_pe_21_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_21),
		.in_col (out_col_20_22),
		.out_row (out_row_21_22),
		.out_col (out_col_21_22),
		.out_data (out_data_21_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_23;
	wire signed [DATA_WIDTH-1:0] out_col_21_23;
	wire signed [DATA_WIDTH-1:0] out_data_21_23;
	integer_mac_pe mac_pe_21_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_22),
		.in_col (out_col_20_23),
		.out_row (out_row_21_23),
		.out_col (out_col_21_23),
		.out_data (out_data_21_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_24;
	wire signed [DATA_WIDTH-1:0] out_col_21_24;
	wire signed [DATA_WIDTH-1:0] out_data_21_24;
	integer_mac_pe mac_pe_21_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_23),
		.in_col (out_col_20_24),
		.out_row (out_row_21_24),
		.out_col (out_col_21_24),
		.out_data (out_data_21_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_25;
	wire signed [DATA_WIDTH-1:0] out_col_21_25;
	wire signed [DATA_WIDTH-1:0] out_data_21_25;
	integer_mac_pe mac_pe_21_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_24),
		.in_col (out_col_20_25),
		.out_row (out_row_21_25),
		.out_col (out_col_21_25),
		.out_data (out_data_21_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_26;
	wire signed [DATA_WIDTH-1:0] out_col_21_26;
	wire signed [DATA_WIDTH-1:0] out_data_21_26;
	integer_mac_pe mac_pe_21_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_25),
		.in_col (out_col_20_26),
		.out_row (out_row_21_26),
		.out_col (out_col_21_26),
		.out_data (out_data_21_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_27;
	wire signed [DATA_WIDTH-1:0] out_col_21_27;
	wire signed [DATA_WIDTH-1:0] out_data_21_27;
	integer_mac_pe mac_pe_21_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_26),
		.in_col (out_col_20_27),
		.out_row (out_row_21_27),
		.out_col (out_col_21_27),
		.out_data (out_data_21_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_28;
	wire signed [DATA_WIDTH-1:0] out_col_21_28;
	wire signed [DATA_WIDTH-1:0] out_data_21_28;
	integer_mac_pe mac_pe_21_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_27),
		.in_col (out_col_20_28),
		.out_row (out_row_21_28),
		.out_col (out_col_21_28),
		.out_data (out_data_21_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_29;
	wire signed [DATA_WIDTH-1:0] out_col_21_29;
	wire signed [DATA_WIDTH-1:0] out_data_21_29;
	integer_mac_pe mac_pe_21_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_28),
		.in_col (out_col_20_29),
		.out_row (out_row_21_29),
		.out_col (out_col_21_29),
		.out_data (out_data_21_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_30;
	wire signed [DATA_WIDTH-1:0] out_col_21_30;
	wire signed [DATA_WIDTH-1:0] out_data_21_30;
	integer_mac_pe mac_pe_21_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_29),
		.in_col (out_col_20_30),
		.out_row (out_row_21_30),
		.out_col (out_col_21_30),
		.out_data (out_data_21_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_21_31;
	wire signed [DATA_WIDTH-1:0] out_col_21_31;
	wire signed [DATA_WIDTH-1:0] out_data_21_31;
	integer_mac_pe mac_pe_21_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_21_30),
		.in_col (out_col_20_31),
		.out_row (out_row_21_31),
		.out_col (out_col_21_31),
		.out_data (out_data_21_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_0;
	wire signed [DATA_WIDTH-1:0] out_col_22_0;
	wire signed [DATA_WIDTH-1:0] out_data_22_0;
	integer_mac_pe mac_pe_22_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_22_out),
		.in_col (out_col_21_0),
		.out_row (out_row_22_0),
		.out_col (out_col_22_0),
		.out_data (out_data_22_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_1;
	wire signed [DATA_WIDTH-1:0] out_col_22_1;
	wire signed [DATA_WIDTH-1:0] out_data_22_1;
	integer_mac_pe mac_pe_22_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_0),
		.in_col (out_col_21_1),
		.out_row (out_row_22_1),
		.out_col (out_col_22_1),
		.out_data (out_data_22_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_2;
	wire signed [DATA_WIDTH-1:0] out_col_22_2;
	wire signed [DATA_WIDTH-1:0] out_data_22_2;
	integer_mac_pe mac_pe_22_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_1),
		.in_col (out_col_21_2),
		.out_row (out_row_22_2),
		.out_col (out_col_22_2),
		.out_data (out_data_22_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_3;
	wire signed [DATA_WIDTH-1:0] out_col_22_3;
	wire signed [DATA_WIDTH-1:0] out_data_22_3;
	integer_mac_pe mac_pe_22_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_2),
		.in_col (out_col_21_3),
		.out_row (out_row_22_3),
		.out_col (out_col_22_3),
		.out_data (out_data_22_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_4;
	wire signed [DATA_WIDTH-1:0] out_col_22_4;
	wire signed [DATA_WIDTH-1:0] out_data_22_4;
	integer_mac_pe mac_pe_22_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_3),
		.in_col (out_col_21_4),
		.out_row (out_row_22_4),
		.out_col (out_col_22_4),
		.out_data (out_data_22_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_5;
	wire signed [DATA_WIDTH-1:0] out_col_22_5;
	wire signed [DATA_WIDTH-1:0] out_data_22_5;
	integer_mac_pe mac_pe_22_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_4),
		.in_col (out_col_21_5),
		.out_row (out_row_22_5),
		.out_col (out_col_22_5),
		.out_data (out_data_22_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_6;
	wire signed [DATA_WIDTH-1:0] out_col_22_6;
	wire signed [DATA_WIDTH-1:0] out_data_22_6;
	integer_mac_pe mac_pe_22_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_5),
		.in_col (out_col_21_6),
		.out_row (out_row_22_6),
		.out_col (out_col_22_6),
		.out_data (out_data_22_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_7;
	wire signed [DATA_WIDTH-1:0] out_col_22_7;
	wire signed [DATA_WIDTH-1:0] out_data_22_7;
	integer_mac_pe mac_pe_22_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_6),
		.in_col (out_col_21_7),
		.out_row (out_row_22_7),
		.out_col (out_col_22_7),
		.out_data (out_data_22_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_8;
	wire signed [DATA_WIDTH-1:0] out_col_22_8;
	wire signed [DATA_WIDTH-1:0] out_data_22_8;
	integer_mac_pe mac_pe_22_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_7),
		.in_col (out_col_21_8),
		.out_row (out_row_22_8),
		.out_col (out_col_22_8),
		.out_data (out_data_22_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_9;
	wire signed [DATA_WIDTH-1:0] out_col_22_9;
	wire signed [DATA_WIDTH-1:0] out_data_22_9;
	integer_mac_pe mac_pe_22_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_8),
		.in_col (out_col_21_9),
		.out_row (out_row_22_9),
		.out_col (out_col_22_9),
		.out_data (out_data_22_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_10;
	wire signed [DATA_WIDTH-1:0] out_col_22_10;
	wire signed [DATA_WIDTH-1:0] out_data_22_10;
	integer_mac_pe mac_pe_22_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_9),
		.in_col (out_col_21_10),
		.out_row (out_row_22_10),
		.out_col (out_col_22_10),
		.out_data (out_data_22_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_11;
	wire signed [DATA_WIDTH-1:0] out_col_22_11;
	wire signed [DATA_WIDTH-1:0] out_data_22_11;
	integer_mac_pe mac_pe_22_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_10),
		.in_col (out_col_21_11),
		.out_row (out_row_22_11),
		.out_col (out_col_22_11),
		.out_data (out_data_22_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_12;
	wire signed [DATA_WIDTH-1:0] out_col_22_12;
	wire signed [DATA_WIDTH-1:0] out_data_22_12;
	integer_mac_pe mac_pe_22_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_11),
		.in_col (out_col_21_12),
		.out_row (out_row_22_12),
		.out_col (out_col_22_12),
		.out_data (out_data_22_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_13;
	wire signed [DATA_WIDTH-1:0] out_col_22_13;
	wire signed [DATA_WIDTH-1:0] out_data_22_13;
	integer_mac_pe mac_pe_22_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_12),
		.in_col (out_col_21_13),
		.out_row (out_row_22_13),
		.out_col (out_col_22_13),
		.out_data (out_data_22_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_14;
	wire signed [DATA_WIDTH-1:0] out_col_22_14;
	wire signed [DATA_WIDTH-1:0] out_data_22_14;
	integer_mac_pe mac_pe_22_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_13),
		.in_col (out_col_21_14),
		.out_row (out_row_22_14),
		.out_col (out_col_22_14),
		.out_data (out_data_22_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_15;
	wire signed [DATA_WIDTH-1:0] out_col_22_15;
	wire signed [DATA_WIDTH-1:0] out_data_22_15;
	integer_mac_pe mac_pe_22_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_14),
		.in_col (out_col_21_15),
		.out_row (out_row_22_15),
		.out_col (out_col_22_15),
		.out_data (out_data_22_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_16;
	wire signed [DATA_WIDTH-1:0] out_col_22_16;
	wire signed [DATA_WIDTH-1:0] out_data_22_16;
	integer_mac_pe mac_pe_22_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_15),
		.in_col (out_col_21_16),
		.out_row (out_row_22_16),
		.out_col (out_col_22_16),
		.out_data (out_data_22_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_17;
	wire signed [DATA_WIDTH-1:0] out_col_22_17;
	wire signed [DATA_WIDTH-1:0] out_data_22_17;
	integer_mac_pe mac_pe_22_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_16),
		.in_col (out_col_21_17),
		.out_row (out_row_22_17),
		.out_col (out_col_22_17),
		.out_data (out_data_22_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_18;
	wire signed [DATA_WIDTH-1:0] out_col_22_18;
	wire signed [DATA_WIDTH-1:0] out_data_22_18;
	integer_mac_pe mac_pe_22_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_17),
		.in_col (out_col_21_18),
		.out_row (out_row_22_18),
		.out_col (out_col_22_18),
		.out_data (out_data_22_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_19;
	wire signed [DATA_WIDTH-1:0] out_col_22_19;
	wire signed [DATA_WIDTH-1:0] out_data_22_19;
	integer_mac_pe mac_pe_22_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_18),
		.in_col (out_col_21_19),
		.out_row (out_row_22_19),
		.out_col (out_col_22_19),
		.out_data (out_data_22_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_20;
	wire signed [DATA_WIDTH-1:0] out_col_22_20;
	wire signed [DATA_WIDTH-1:0] out_data_22_20;
	integer_mac_pe mac_pe_22_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_19),
		.in_col (out_col_21_20),
		.out_row (out_row_22_20),
		.out_col (out_col_22_20),
		.out_data (out_data_22_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_21;
	wire signed [DATA_WIDTH-1:0] out_col_22_21;
	wire signed [DATA_WIDTH-1:0] out_data_22_21;
	integer_mac_pe mac_pe_22_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_20),
		.in_col (out_col_21_21),
		.out_row (out_row_22_21),
		.out_col (out_col_22_21),
		.out_data (out_data_22_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_22;
	wire signed [DATA_WIDTH-1:0] out_col_22_22;
	wire signed [DATA_WIDTH-1:0] out_data_22_22;
	integer_mac_pe mac_pe_22_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_21),
		.in_col (out_col_21_22),
		.out_row (out_row_22_22),
		.out_col (out_col_22_22),
		.out_data (out_data_22_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_23;
	wire signed [DATA_WIDTH-1:0] out_col_22_23;
	wire signed [DATA_WIDTH-1:0] out_data_22_23;
	integer_mac_pe mac_pe_22_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_22),
		.in_col (out_col_21_23),
		.out_row (out_row_22_23),
		.out_col (out_col_22_23),
		.out_data (out_data_22_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_24;
	wire signed [DATA_WIDTH-1:0] out_col_22_24;
	wire signed [DATA_WIDTH-1:0] out_data_22_24;
	integer_mac_pe mac_pe_22_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_23),
		.in_col (out_col_21_24),
		.out_row (out_row_22_24),
		.out_col (out_col_22_24),
		.out_data (out_data_22_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_25;
	wire signed [DATA_WIDTH-1:0] out_col_22_25;
	wire signed [DATA_WIDTH-1:0] out_data_22_25;
	integer_mac_pe mac_pe_22_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_24),
		.in_col (out_col_21_25),
		.out_row (out_row_22_25),
		.out_col (out_col_22_25),
		.out_data (out_data_22_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_26;
	wire signed [DATA_WIDTH-1:0] out_col_22_26;
	wire signed [DATA_WIDTH-1:0] out_data_22_26;
	integer_mac_pe mac_pe_22_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_25),
		.in_col (out_col_21_26),
		.out_row (out_row_22_26),
		.out_col (out_col_22_26),
		.out_data (out_data_22_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_27;
	wire signed [DATA_WIDTH-1:0] out_col_22_27;
	wire signed [DATA_WIDTH-1:0] out_data_22_27;
	integer_mac_pe mac_pe_22_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_26),
		.in_col (out_col_21_27),
		.out_row (out_row_22_27),
		.out_col (out_col_22_27),
		.out_data (out_data_22_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_28;
	wire signed [DATA_WIDTH-1:0] out_col_22_28;
	wire signed [DATA_WIDTH-1:0] out_data_22_28;
	integer_mac_pe mac_pe_22_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_27),
		.in_col (out_col_21_28),
		.out_row (out_row_22_28),
		.out_col (out_col_22_28),
		.out_data (out_data_22_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_29;
	wire signed [DATA_WIDTH-1:0] out_col_22_29;
	wire signed [DATA_WIDTH-1:0] out_data_22_29;
	integer_mac_pe mac_pe_22_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_28),
		.in_col (out_col_21_29),
		.out_row (out_row_22_29),
		.out_col (out_col_22_29),
		.out_data (out_data_22_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_30;
	wire signed [DATA_WIDTH-1:0] out_col_22_30;
	wire signed [DATA_WIDTH-1:0] out_data_22_30;
	integer_mac_pe mac_pe_22_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_29),
		.in_col (out_col_21_30),
		.out_row (out_row_22_30),
		.out_col (out_col_22_30),
		.out_data (out_data_22_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_22_31;
	wire signed [DATA_WIDTH-1:0] out_col_22_31;
	wire signed [DATA_WIDTH-1:0] out_data_22_31;
	integer_mac_pe mac_pe_22_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_22_30),
		.in_col (out_col_21_31),
		.out_row (out_row_22_31),
		.out_col (out_col_22_31),
		.out_data (out_data_22_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_0;
	wire signed [DATA_WIDTH-1:0] out_col_23_0;
	wire signed [DATA_WIDTH-1:0] out_data_23_0;
	integer_mac_pe mac_pe_23_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_23_out),
		.in_col (out_col_22_0),
		.out_row (out_row_23_0),
		.out_col (out_col_23_0),
		.out_data (out_data_23_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_1;
	wire signed [DATA_WIDTH-1:0] out_col_23_1;
	wire signed [DATA_WIDTH-1:0] out_data_23_1;
	integer_mac_pe mac_pe_23_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_0),
		.in_col (out_col_22_1),
		.out_row (out_row_23_1),
		.out_col (out_col_23_1),
		.out_data (out_data_23_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_2;
	wire signed [DATA_WIDTH-1:0] out_col_23_2;
	wire signed [DATA_WIDTH-1:0] out_data_23_2;
	integer_mac_pe mac_pe_23_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_1),
		.in_col (out_col_22_2),
		.out_row (out_row_23_2),
		.out_col (out_col_23_2),
		.out_data (out_data_23_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_3;
	wire signed [DATA_WIDTH-1:0] out_col_23_3;
	wire signed [DATA_WIDTH-1:0] out_data_23_3;
	integer_mac_pe mac_pe_23_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_2),
		.in_col (out_col_22_3),
		.out_row (out_row_23_3),
		.out_col (out_col_23_3),
		.out_data (out_data_23_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_4;
	wire signed [DATA_WIDTH-1:0] out_col_23_4;
	wire signed [DATA_WIDTH-1:0] out_data_23_4;
	integer_mac_pe mac_pe_23_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_3),
		.in_col (out_col_22_4),
		.out_row (out_row_23_4),
		.out_col (out_col_23_4),
		.out_data (out_data_23_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_5;
	wire signed [DATA_WIDTH-1:0] out_col_23_5;
	wire signed [DATA_WIDTH-1:0] out_data_23_5;
	integer_mac_pe mac_pe_23_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_4),
		.in_col (out_col_22_5),
		.out_row (out_row_23_5),
		.out_col (out_col_23_5),
		.out_data (out_data_23_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_6;
	wire signed [DATA_WIDTH-1:0] out_col_23_6;
	wire signed [DATA_WIDTH-1:0] out_data_23_6;
	integer_mac_pe mac_pe_23_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_5),
		.in_col (out_col_22_6),
		.out_row (out_row_23_6),
		.out_col (out_col_23_6),
		.out_data (out_data_23_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_7;
	wire signed [DATA_WIDTH-1:0] out_col_23_7;
	wire signed [DATA_WIDTH-1:0] out_data_23_7;
	integer_mac_pe mac_pe_23_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_6),
		.in_col (out_col_22_7),
		.out_row (out_row_23_7),
		.out_col (out_col_23_7),
		.out_data (out_data_23_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_8;
	wire signed [DATA_WIDTH-1:0] out_col_23_8;
	wire signed [DATA_WIDTH-1:0] out_data_23_8;
	integer_mac_pe mac_pe_23_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_7),
		.in_col (out_col_22_8),
		.out_row (out_row_23_8),
		.out_col (out_col_23_8),
		.out_data (out_data_23_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_9;
	wire signed [DATA_WIDTH-1:0] out_col_23_9;
	wire signed [DATA_WIDTH-1:0] out_data_23_9;
	integer_mac_pe mac_pe_23_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_8),
		.in_col (out_col_22_9),
		.out_row (out_row_23_9),
		.out_col (out_col_23_9),
		.out_data (out_data_23_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_10;
	wire signed [DATA_WIDTH-1:0] out_col_23_10;
	wire signed [DATA_WIDTH-1:0] out_data_23_10;
	integer_mac_pe mac_pe_23_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_9),
		.in_col (out_col_22_10),
		.out_row (out_row_23_10),
		.out_col (out_col_23_10),
		.out_data (out_data_23_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_11;
	wire signed [DATA_WIDTH-1:0] out_col_23_11;
	wire signed [DATA_WIDTH-1:0] out_data_23_11;
	integer_mac_pe mac_pe_23_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_10),
		.in_col (out_col_22_11),
		.out_row (out_row_23_11),
		.out_col (out_col_23_11),
		.out_data (out_data_23_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_12;
	wire signed [DATA_WIDTH-1:0] out_col_23_12;
	wire signed [DATA_WIDTH-1:0] out_data_23_12;
	integer_mac_pe mac_pe_23_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_11),
		.in_col (out_col_22_12),
		.out_row (out_row_23_12),
		.out_col (out_col_23_12),
		.out_data (out_data_23_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_13;
	wire signed [DATA_WIDTH-1:0] out_col_23_13;
	wire signed [DATA_WIDTH-1:0] out_data_23_13;
	integer_mac_pe mac_pe_23_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_12),
		.in_col (out_col_22_13),
		.out_row (out_row_23_13),
		.out_col (out_col_23_13),
		.out_data (out_data_23_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_14;
	wire signed [DATA_WIDTH-1:0] out_col_23_14;
	wire signed [DATA_WIDTH-1:0] out_data_23_14;
	integer_mac_pe mac_pe_23_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_13),
		.in_col (out_col_22_14),
		.out_row (out_row_23_14),
		.out_col (out_col_23_14),
		.out_data (out_data_23_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_15;
	wire signed [DATA_WIDTH-1:0] out_col_23_15;
	wire signed [DATA_WIDTH-1:0] out_data_23_15;
	integer_mac_pe mac_pe_23_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_14),
		.in_col (out_col_22_15),
		.out_row (out_row_23_15),
		.out_col (out_col_23_15),
		.out_data (out_data_23_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_16;
	wire signed [DATA_WIDTH-1:0] out_col_23_16;
	wire signed [DATA_WIDTH-1:0] out_data_23_16;
	integer_mac_pe mac_pe_23_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_15),
		.in_col (out_col_22_16),
		.out_row (out_row_23_16),
		.out_col (out_col_23_16),
		.out_data (out_data_23_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_17;
	wire signed [DATA_WIDTH-1:0] out_col_23_17;
	wire signed [DATA_WIDTH-1:0] out_data_23_17;
	integer_mac_pe mac_pe_23_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_16),
		.in_col (out_col_22_17),
		.out_row (out_row_23_17),
		.out_col (out_col_23_17),
		.out_data (out_data_23_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_18;
	wire signed [DATA_WIDTH-1:0] out_col_23_18;
	wire signed [DATA_WIDTH-1:0] out_data_23_18;
	integer_mac_pe mac_pe_23_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_17),
		.in_col (out_col_22_18),
		.out_row (out_row_23_18),
		.out_col (out_col_23_18),
		.out_data (out_data_23_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_19;
	wire signed [DATA_WIDTH-1:0] out_col_23_19;
	wire signed [DATA_WIDTH-1:0] out_data_23_19;
	integer_mac_pe mac_pe_23_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_18),
		.in_col (out_col_22_19),
		.out_row (out_row_23_19),
		.out_col (out_col_23_19),
		.out_data (out_data_23_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_20;
	wire signed [DATA_WIDTH-1:0] out_col_23_20;
	wire signed [DATA_WIDTH-1:0] out_data_23_20;
	integer_mac_pe mac_pe_23_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_19),
		.in_col (out_col_22_20),
		.out_row (out_row_23_20),
		.out_col (out_col_23_20),
		.out_data (out_data_23_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_21;
	wire signed [DATA_WIDTH-1:0] out_col_23_21;
	wire signed [DATA_WIDTH-1:0] out_data_23_21;
	integer_mac_pe mac_pe_23_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_20),
		.in_col (out_col_22_21),
		.out_row (out_row_23_21),
		.out_col (out_col_23_21),
		.out_data (out_data_23_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_22;
	wire signed [DATA_WIDTH-1:0] out_col_23_22;
	wire signed [DATA_WIDTH-1:0] out_data_23_22;
	integer_mac_pe mac_pe_23_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_21),
		.in_col (out_col_22_22),
		.out_row (out_row_23_22),
		.out_col (out_col_23_22),
		.out_data (out_data_23_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_23;
	wire signed [DATA_WIDTH-1:0] out_col_23_23;
	wire signed [DATA_WIDTH-1:0] out_data_23_23;
	integer_mac_pe mac_pe_23_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_22),
		.in_col (out_col_22_23),
		.out_row (out_row_23_23),
		.out_col (out_col_23_23),
		.out_data (out_data_23_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_24;
	wire signed [DATA_WIDTH-1:0] out_col_23_24;
	wire signed [DATA_WIDTH-1:0] out_data_23_24;
	integer_mac_pe mac_pe_23_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_23),
		.in_col (out_col_22_24),
		.out_row (out_row_23_24),
		.out_col (out_col_23_24),
		.out_data (out_data_23_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_25;
	wire signed [DATA_WIDTH-1:0] out_col_23_25;
	wire signed [DATA_WIDTH-1:0] out_data_23_25;
	integer_mac_pe mac_pe_23_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_24),
		.in_col (out_col_22_25),
		.out_row (out_row_23_25),
		.out_col (out_col_23_25),
		.out_data (out_data_23_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_26;
	wire signed [DATA_WIDTH-1:0] out_col_23_26;
	wire signed [DATA_WIDTH-1:0] out_data_23_26;
	integer_mac_pe mac_pe_23_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_25),
		.in_col (out_col_22_26),
		.out_row (out_row_23_26),
		.out_col (out_col_23_26),
		.out_data (out_data_23_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_27;
	wire signed [DATA_WIDTH-1:0] out_col_23_27;
	wire signed [DATA_WIDTH-1:0] out_data_23_27;
	integer_mac_pe mac_pe_23_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_26),
		.in_col (out_col_22_27),
		.out_row (out_row_23_27),
		.out_col (out_col_23_27),
		.out_data (out_data_23_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_28;
	wire signed [DATA_WIDTH-1:0] out_col_23_28;
	wire signed [DATA_WIDTH-1:0] out_data_23_28;
	integer_mac_pe mac_pe_23_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_27),
		.in_col (out_col_22_28),
		.out_row (out_row_23_28),
		.out_col (out_col_23_28),
		.out_data (out_data_23_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_29;
	wire signed [DATA_WIDTH-1:0] out_col_23_29;
	wire signed [DATA_WIDTH-1:0] out_data_23_29;
	integer_mac_pe mac_pe_23_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_28),
		.in_col (out_col_22_29),
		.out_row (out_row_23_29),
		.out_col (out_col_23_29),
		.out_data (out_data_23_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_30;
	wire signed [DATA_WIDTH-1:0] out_col_23_30;
	wire signed [DATA_WIDTH-1:0] out_data_23_30;
	integer_mac_pe mac_pe_23_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_29),
		.in_col (out_col_22_30),
		.out_row (out_row_23_30),
		.out_col (out_col_23_30),
		.out_data (out_data_23_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_23_31;
	wire signed [DATA_WIDTH-1:0] out_col_23_31;
	wire signed [DATA_WIDTH-1:0] out_data_23_31;
	integer_mac_pe mac_pe_23_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_23_30),
		.in_col (out_col_22_31),
		.out_row (out_row_23_31),
		.out_col (out_col_23_31),
		.out_data (out_data_23_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_0;
	wire signed [DATA_WIDTH-1:0] out_col_24_0;
	wire signed [DATA_WIDTH-1:0] out_data_24_0;
	integer_mac_pe mac_pe_24_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_24_out),
		.in_col (out_col_23_0),
		.out_row (out_row_24_0),
		.out_col (out_col_24_0),
		.out_data (out_data_24_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_1;
	wire signed [DATA_WIDTH-1:0] out_col_24_1;
	wire signed [DATA_WIDTH-1:0] out_data_24_1;
	integer_mac_pe mac_pe_24_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_0),
		.in_col (out_col_23_1),
		.out_row (out_row_24_1),
		.out_col (out_col_24_1),
		.out_data (out_data_24_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_2;
	wire signed [DATA_WIDTH-1:0] out_col_24_2;
	wire signed [DATA_WIDTH-1:0] out_data_24_2;
	integer_mac_pe mac_pe_24_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_1),
		.in_col (out_col_23_2),
		.out_row (out_row_24_2),
		.out_col (out_col_24_2),
		.out_data (out_data_24_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_3;
	wire signed [DATA_WIDTH-1:0] out_col_24_3;
	wire signed [DATA_WIDTH-1:0] out_data_24_3;
	integer_mac_pe mac_pe_24_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_2),
		.in_col (out_col_23_3),
		.out_row (out_row_24_3),
		.out_col (out_col_24_3),
		.out_data (out_data_24_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_4;
	wire signed [DATA_WIDTH-1:0] out_col_24_4;
	wire signed [DATA_WIDTH-1:0] out_data_24_4;
	integer_mac_pe mac_pe_24_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_3),
		.in_col (out_col_23_4),
		.out_row (out_row_24_4),
		.out_col (out_col_24_4),
		.out_data (out_data_24_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_5;
	wire signed [DATA_WIDTH-1:0] out_col_24_5;
	wire signed [DATA_WIDTH-1:0] out_data_24_5;
	integer_mac_pe mac_pe_24_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_4),
		.in_col (out_col_23_5),
		.out_row (out_row_24_5),
		.out_col (out_col_24_5),
		.out_data (out_data_24_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_6;
	wire signed [DATA_WIDTH-1:0] out_col_24_6;
	wire signed [DATA_WIDTH-1:0] out_data_24_6;
	integer_mac_pe mac_pe_24_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_5),
		.in_col (out_col_23_6),
		.out_row (out_row_24_6),
		.out_col (out_col_24_6),
		.out_data (out_data_24_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_7;
	wire signed [DATA_WIDTH-1:0] out_col_24_7;
	wire signed [DATA_WIDTH-1:0] out_data_24_7;
	integer_mac_pe mac_pe_24_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_6),
		.in_col (out_col_23_7),
		.out_row (out_row_24_7),
		.out_col (out_col_24_7),
		.out_data (out_data_24_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_8;
	wire signed [DATA_WIDTH-1:0] out_col_24_8;
	wire signed [DATA_WIDTH-1:0] out_data_24_8;
	integer_mac_pe mac_pe_24_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_7),
		.in_col (out_col_23_8),
		.out_row (out_row_24_8),
		.out_col (out_col_24_8),
		.out_data (out_data_24_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_9;
	wire signed [DATA_WIDTH-1:0] out_col_24_9;
	wire signed [DATA_WIDTH-1:0] out_data_24_9;
	integer_mac_pe mac_pe_24_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_8),
		.in_col (out_col_23_9),
		.out_row (out_row_24_9),
		.out_col (out_col_24_9),
		.out_data (out_data_24_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_10;
	wire signed [DATA_WIDTH-1:0] out_col_24_10;
	wire signed [DATA_WIDTH-1:0] out_data_24_10;
	integer_mac_pe mac_pe_24_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_9),
		.in_col (out_col_23_10),
		.out_row (out_row_24_10),
		.out_col (out_col_24_10),
		.out_data (out_data_24_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_11;
	wire signed [DATA_WIDTH-1:0] out_col_24_11;
	wire signed [DATA_WIDTH-1:0] out_data_24_11;
	integer_mac_pe mac_pe_24_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_10),
		.in_col (out_col_23_11),
		.out_row (out_row_24_11),
		.out_col (out_col_24_11),
		.out_data (out_data_24_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_12;
	wire signed [DATA_WIDTH-1:0] out_col_24_12;
	wire signed [DATA_WIDTH-1:0] out_data_24_12;
	integer_mac_pe mac_pe_24_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_11),
		.in_col (out_col_23_12),
		.out_row (out_row_24_12),
		.out_col (out_col_24_12),
		.out_data (out_data_24_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_13;
	wire signed [DATA_WIDTH-1:0] out_col_24_13;
	wire signed [DATA_WIDTH-1:0] out_data_24_13;
	integer_mac_pe mac_pe_24_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_12),
		.in_col (out_col_23_13),
		.out_row (out_row_24_13),
		.out_col (out_col_24_13),
		.out_data (out_data_24_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_14;
	wire signed [DATA_WIDTH-1:0] out_col_24_14;
	wire signed [DATA_WIDTH-1:0] out_data_24_14;
	integer_mac_pe mac_pe_24_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_13),
		.in_col (out_col_23_14),
		.out_row (out_row_24_14),
		.out_col (out_col_24_14),
		.out_data (out_data_24_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_15;
	wire signed [DATA_WIDTH-1:0] out_col_24_15;
	wire signed [DATA_WIDTH-1:0] out_data_24_15;
	integer_mac_pe mac_pe_24_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_14),
		.in_col (out_col_23_15),
		.out_row (out_row_24_15),
		.out_col (out_col_24_15),
		.out_data (out_data_24_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_16;
	wire signed [DATA_WIDTH-1:0] out_col_24_16;
	wire signed [DATA_WIDTH-1:0] out_data_24_16;
	integer_mac_pe mac_pe_24_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_15),
		.in_col (out_col_23_16),
		.out_row (out_row_24_16),
		.out_col (out_col_24_16),
		.out_data (out_data_24_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_17;
	wire signed [DATA_WIDTH-1:0] out_col_24_17;
	wire signed [DATA_WIDTH-1:0] out_data_24_17;
	integer_mac_pe mac_pe_24_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_16),
		.in_col (out_col_23_17),
		.out_row (out_row_24_17),
		.out_col (out_col_24_17),
		.out_data (out_data_24_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_18;
	wire signed [DATA_WIDTH-1:0] out_col_24_18;
	wire signed [DATA_WIDTH-1:0] out_data_24_18;
	integer_mac_pe mac_pe_24_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_17),
		.in_col (out_col_23_18),
		.out_row (out_row_24_18),
		.out_col (out_col_24_18),
		.out_data (out_data_24_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_19;
	wire signed [DATA_WIDTH-1:0] out_col_24_19;
	wire signed [DATA_WIDTH-1:0] out_data_24_19;
	integer_mac_pe mac_pe_24_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_18),
		.in_col (out_col_23_19),
		.out_row (out_row_24_19),
		.out_col (out_col_24_19),
		.out_data (out_data_24_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_20;
	wire signed [DATA_WIDTH-1:0] out_col_24_20;
	wire signed [DATA_WIDTH-1:0] out_data_24_20;
	integer_mac_pe mac_pe_24_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_19),
		.in_col (out_col_23_20),
		.out_row (out_row_24_20),
		.out_col (out_col_24_20),
		.out_data (out_data_24_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_21;
	wire signed [DATA_WIDTH-1:0] out_col_24_21;
	wire signed [DATA_WIDTH-1:0] out_data_24_21;
	integer_mac_pe mac_pe_24_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_20),
		.in_col (out_col_23_21),
		.out_row (out_row_24_21),
		.out_col (out_col_24_21),
		.out_data (out_data_24_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_22;
	wire signed [DATA_WIDTH-1:0] out_col_24_22;
	wire signed [DATA_WIDTH-1:0] out_data_24_22;
	integer_mac_pe mac_pe_24_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_21),
		.in_col (out_col_23_22),
		.out_row (out_row_24_22),
		.out_col (out_col_24_22),
		.out_data (out_data_24_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_23;
	wire signed [DATA_WIDTH-1:0] out_col_24_23;
	wire signed [DATA_WIDTH-1:0] out_data_24_23;
	integer_mac_pe mac_pe_24_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_22),
		.in_col (out_col_23_23),
		.out_row (out_row_24_23),
		.out_col (out_col_24_23),
		.out_data (out_data_24_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_24;
	wire signed [DATA_WIDTH-1:0] out_col_24_24;
	wire signed [DATA_WIDTH-1:0] out_data_24_24;
	integer_mac_pe mac_pe_24_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_23),
		.in_col (out_col_23_24),
		.out_row (out_row_24_24),
		.out_col (out_col_24_24),
		.out_data (out_data_24_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_25;
	wire signed [DATA_WIDTH-1:0] out_col_24_25;
	wire signed [DATA_WIDTH-1:0] out_data_24_25;
	integer_mac_pe mac_pe_24_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_24),
		.in_col (out_col_23_25),
		.out_row (out_row_24_25),
		.out_col (out_col_24_25),
		.out_data (out_data_24_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_26;
	wire signed [DATA_WIDTH-1:0] out_col_24_26;
	wire signed [DATA_WIDTH-1:0] out_data_24_26;
	integer_mac_pe mac_pe_24_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_25),
		.in_col (out_col_23_26),
		.out_row (out_row_24_26),
		.out_col (out_col_24_26),
		.out_data (out_data_24_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_27;
	wire signed [DATA_WIDTH-1:0] out_col_24_27;
	wire signed [DATA_WIDTH-1:0] out_data_24_27;
	integer_mac_pe mac_pe_24_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_26),
		.in_col (out_col_23_27),
		.out_row (out_row_24_27),
		.out_col (out_col_24_27),
		.out_data (out_data_24_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_28;
	wire signed [DATA_WIDTH-1:0] out_col_24_28;
	wire signed [DATA_WIDTH-1:0] out_data_24_28;
	integer_mac_pe mac_pe_24_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_27),
		.in_col (out_col_23_28),
		.out_row (out_row_24_28),
		.out_col (out_col_24_28),
		.out_data (out_data_24_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_29;
	wire signed [DATA_WIDTH-1:0] out_col_24_29;
	wire signed [DATA_WIDTH-1:0] out_data_24_29;
	integer_mac_pe mac_pe_24_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_28),
		.in_col (out_col_23_29),
		.out_row (out_row_24_29),
		.out_col (out_col_24_29),
		.out_data (out_data_24_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_30;
	wire signed [DATA_WIDTH-1:0] out_col_24_30;
	wire signed [DATA_WIDTH-1:0] out_data_24_30;
	integer_mac_pe mac_pe_24_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_29),
		.in_col (out_col_23_30),
		.out_row (out_row_24_30),
		.out_col (out_col_24_30),
		.out_data (out_data_24_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_24_31;
	wire signed [DATA_WIDTH-1:0] out_col_24_31;
	wire signed [DATA_WIDTH-1:0] out_data_24_31;
	integer_mac_pe mac_pe_24_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_24_30),
		.in_col (out_col_23_31),
		.out_row (out_row_24_31),
		.out_col (out_col_24_31),
		.out_data (out_data_24_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_0;
	wire signed [DATA_WIDTH-1:0] out_col_25_0;
	wire signed [DATA_WIDTH-1:0] out_data_25_0;
	integer_mac_pe mac_pe_25_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_25_out),
		.in_col (out_col_24_0),
		.out_row (out_row_25_0),
		.out_col (out_col_25_0),
		.out_data (out_data_25_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_1;
	wire signed [DATA_WIDTH-1:0] out_col_25_1;
	wire signed [DATA_WIDTH-1:0] out_data_25_1;
	integer_mac_pe mac_pe_25_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_0),
		.in_col (out_col_24_1),
		.out_row (out_row_25_1),
		.out_col (out_col_25_1),
		.out_data (out_data_25_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_2;
	wire signed [DATA_WIDTH-1:0] out_col_25_2;
	wire signed [DATA_WIDTH-1:0] out_data_25_2;
	integer_mac_pe mac_pe_25_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_1),
		.in_col (out_col_24_2),
		.out_row (out_row_25_2),
		.out_col (out_col_25_2),
		.out_data (out_data_25_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_3;
	wire signed [DATA_WIDTH-1:0] out_col_25_3;
	wire signed [DATA_WIDTH-1:0] out_data_25_3;
	integer_mac_pe mac_pe_25_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_2),
		.in_col (out_col_24_3),
		.out_row (out_row_25_3),
		.out_col (out_col_25_3),
		.out_data (out_data_25_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_4;
	wire signed [DATA_WIDTH-1:0] out_col_25_4;
	wire signed [DATA_WIDTH-1:0] out_data_25_4;
	integer_mac_pe mac_pe_25_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_3),
		.in_col (out_col_24_4),
		.out_row (out_row_25_4),
		.out_col (out_col_25_4),
		.out_data (out_data_25_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_5;
	wire signed [DATA_WIDTH-1:0] out_col_25_5;
	wire signed [DATA_WIDTH-1:0] out_data_25_5;
	integer_mac_pe mac_pe_25_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_4),
		.in_col (out_col_24_5),
		.out_row (out_row_25_5),
		.out_col (out_col_25_5),
		.out_data (out_data_25_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_6;
	wire signed [DATA_WIDTH-1:0] out_col_25_6;
	wire signed [DATA_WIDTH-1:0] out_data_25_6;
	integer_mac_pe mac_pe_25_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_5),
		.in_col (out_col_24_6),
		.out_row (out_row_25_6),
		.out_col (out_col_25_6),
		.out_data (out_data_25_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_7;
	wire signed [DATA_WIDTH-1:0] out_col_25_7;
	wire signed [DATA_WIDTH-1:0] out_data_25_7;
	integer_mac_pe mac_pe_25_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_6),
		.in_col (out_col_24_7),
		.out_row (out_row_25_7),
		.out_col (out_col_25_7),
		.out_data (out_data_25_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_8;
	wire signed [DATA_WIDTH-1:0] out_col_25_8;
	wire signed [DATA_WIDTH-1:0] out_data_25_8;
	integer_mac_pe mac_pe_25_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_7),
		.in_col (out_col_24_8),
		.out_row (out_row_25_8),
		.out_col (out_col_25_8),
		.out_data (out_data_25_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_9;
	wire signed [DATA_WIDTH-1:0] out_col_25_9;
	wire signed [DATA_WIDTH-1:0] out_data_25_9;
	integer_mac_pe mac_pe_25_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_8),
		.in_col (out_col_24_9),
		.out_row (out_row_25_9),
		.out_col (out_col_25_9),
		.out_data (out_data_25_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_10;
	wire signed [DATA_WIDTH-1:0] out_col_25_10;
	wire signed [DATA_WIDTH-1:0] out_data_25_10;
	integer_mac_pe mac_pe_25_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_9),
		.in_col (out_col_24_10),
		.out_row (out_row_25_10),
		.out_col (out_col_25_10),
		.out_data (out_data_25_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_11;
	wire signed [DATA_WIDTH-1:0] out_col_25_11;
	wire signed [DATA_WIDTH-1:0] out_data_25_11;
	integer_mac_pe mac_pe_25_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_10),
		.in_col (out_col_24_11),
		.out_row (out_row_25_11),
		.out_col (out_col_25_11),
		.out_data (out_data_25_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_12;
	wire signed [DATA_WIDTH-1:0] out_col_25_12;
	wire signed [DATA_WIDTH-1:0] out_data_25_12;
	integer_mac_pe mac_pe_25_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_11),
		.in_col (out_col_24_12),
		.out_row (out_row_25_12),
		.out_col (out_col_25_12),
		.out_data (out_data_25_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_13;
	wire signed [DATA_WIDTH-1:0] out_col_25_13;
	wire signed [DATA_WIDTH-1:0] out_data_25_13;
	integer_mac_pe mac_pe_25_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_12),
		.in_col (out_col_24_13),
		.out_row (out_row_25_13),
		.out_col (out_col_25_13),
		.out_data (out_data_25_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_14;
	wire signed [DATA_WIDTH-1:0] out_col_25_14;
	wire signed [DATA_WIDTH-1:0] out_data_25_14;
	integer_mac_pe mac_pe_25_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_13),
		.in_col (out_col_24_14),
		.out_row (out_row_25_14),
		.out_col (out_col_25_14),
		.out_data (out_data_25_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_15;
	wire signed [DATA_WIDTH-1:0] out_col_25_15;
	wire signed [DATA_WIDTH-1:0] out_data_25_15;
	integer_mac_pe mac_pe_25_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_14),
		.in_col (out_col_24_15),
		.out_row (out_row_25_15),
		.out_col (out_col_25_15),
		.out_data (out_data_25_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_16;
	wire signed [DATA_WIDTH-1:0] out_col_25_16;
	wire signed [DATA_WIDTH-1:0] out_data_25_16;
	integer_mac_pe mac_pe_25_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_15),
		.in_col (out_col_24_16),
		.out_row (out_row_25_16),
		.out_col (out_col_25_16),
		.out_data (out_data_25_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_17;
	wire signed [DATA_WIDTH-1:0] out_col_25_17;
	wire signed [DATA_WIDTH-1:0] out_data_25_17;
	integer_mac_pe mac_pe_25_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_16),
		.in_col (out_col_24_17),
		.out_row (out_row_25_17),
		.out_col (out_col_25_17),
		.out_data (out_data_25_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_18;
	wire signed [DATA_WIDTH-1:0] out_col_25_18;
	wire signed [DATA_WIDTH-1:0] out_data_25_18;
	integer_mac_pe mac_pe_25_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_17),
		.in_col (out_col_24_18),
		.out_row (out_row_25_18),
		.out_col (out_col_25_18),
		.out_data (out_data_25_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_19;
	wire signed [DATA_WIDTH-1:0] out_col_25_19;
	wire signed [DATA_WIDTH-1:0] out_data_25_19;
	integer_mac_pe mac_pe_25_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_18),
		.in_col (out_col_24_19),
		.out_row (out_row_25_19),
		.out_col (out_col_25_19),
		.out_data (out_data_25_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_20;
	wire signed [DATA_WIDTH-1:0] out_col_25_20;
	wire signed [DATA_WIDTH-1:0] out_data_25_20;
	integer_mac_pe mac_pe_25_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_19),
		.in_col (out_col_24_20),
		.out_row (out_row_25_20),
		.out_col (out_col_25_20),
		.out_data (out_data_25_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_21;
	wire signed [DATA_WIDTH-1:0] out_col_25_21;
	wire signed [DATA_WIDTH-1:0] out_data_25_21;
	integer_mac_pe mac_pe_25_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_20),
		.in_col (out_col_24_21),
		.out_row (out_row_25_21),
		.out_col (out_col_25_21),
		.out_data (out_data_25_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_22;
	wire signed [DATA_WIDTH-1:0] out_col_25_22;
	wire signed [DATA_WIDTH-1:0] out_data_25_22;
	integer_mac_pe mac_pe_25_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_21),
		.in_col (out_col_24_22),
		.out_row (out_row_25_22),
		.out_col (out_col_25_22),
		.out_data (out_data_25_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_23;
	wire signed [DATA_WIDTH-1:0] out_col_25_23;
	wire signed [DATA_WIDTH-1:0] out_data_25_23;
	integer_mac_pe mac_pe_25_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_22),
		.in_col (out_col_24_23),
		.out_row (out_row_25_23),
		.out_col (out_col_25_23),
		.out_data (out_data_25_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_24;
	wire signed [DATA_WIDTH-1:0] out_col_25_24;
	wire signed [DATA_WIDTH-1:0] out_data_25_24;
	integer_mac_pe mac_pe_25_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_23),
		.in_col (out_col_24_24),
		.out_row (out_row_25_24),
		.out_col (out_col_25_24),
		.out_data (out_data_25_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_25;
	wire signed [DATA_WIDTH-1:0] out_col_25_25;
	wire signed [DATA_WIDTH-1:0] out_data_25_25;
	integer_mac_pe mac_pe_25_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_24),
		.in_col (out_col_24_25),
		.out_row (out_row_25_25),
		.out_col (out_col_25_25),
		.out_data (out_data_25_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_26;
	wire signed [DATA_WIDTH-1:0] out_col_25_26;
	wire signed [DATA_WIDTH-1:0] out_data_25_26;
	integer_mac_pe mac_pe_25_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_25),
		.in_col (out_col_24_26),
		.out_row (out_row_25_26),
		.out_col (out_col_25_26),
		.out_data (out_data_25_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_27;
	wire signed [DATA_WIDTH-1:0] out_col_25_27;
	wire signed [DATA_WIDTH-1:0] out_data_25_27;
	integer_mac_pe mac_pe_25_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_26),
		.in_col (out_col_24_27),
		.out_row (out_row_25_27),
		.out_col (out_col_25_27),
		.out_data (out_data_25_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_28;
	wire signed [DATA_WIDTH-1:0] out_col_25_28;
	wire signed [DATA_WIDTH-1:0] out_data_25_28;
	integer_mac_pe mac_pe_25_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_27),
		.in_col (out_col_24_28),
		.out_row (out_row_25_28),
		.out_col (out_col_25_28),
		.out_data (out_data_25_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_29;
	wire signed [DATA_WIDTH-1:0] out_col_25_29;
	wire signed [DATA_WIDTH-1:0] out_data_25_29;
	integer_mac_pe mac_pe_25_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_28),
		.in_col (out_col_24_29),
		.out_row (out_row_25_29),
		.out_col (out_col_25_29),
		.out_data (out_data_25_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_30;
	wire signed [DATA_WIDTH-1:0] out_col_25_30;
	wire signed [DATA_WIDTH-1:0] out_data_25_30;
	integer_mac_pe mac_pe_25_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_29),
		.in_col (out_col_24_30),
		.out_row (out_row_25_30),
		.out_col (out_col_25_30),
		.out_data (out_data_25_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_25_31;
	wire signed [DATA_WIDTH-1:0] out_col_25_31;
	wire signed [DATA_WIDTH-1:0] out_data_25_31;
	integer_mac_pe mac_pe_25_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_25_30),
		.in_col (out_col_24_31),
		.out_row (out_row_25_31),
		.out_col (out_col_25_31),
		.out_data (out_data_25_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_0;
	wire signed [DATA_WIDTH-1:0] out_col_26_0;
	wire signed [DATA_WIDTH-1:0] out_data_26_0;
	integer_mac_pe mac_pe_26_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_26_out),
		.in_col (out_col_25_0),
		.out_row (out_row_26_0),
		.out_col (out_col_26_0),
		.out_data (out_data_26_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_1;
	wire signed [DATA_WIDTH-1:0] out_col_26_1;
	wire signed [DATA_WIDTH-1:0] out_data_26_1;
	integer_mac_pe mac_pe_26_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_0),
		.in_col (out_col_25_1),
		.out_row (out_row_26_1),
		.out_col (out_col_26_1),
		.out_data (out_data_26_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_2;
	wire signed [DATA_WIDTH-1:0] out_col_26_2;
	wire signed [DATA_WIDTH-1:0] out_data_26_2;
	integer_mac_pe mac_pe_26_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_1),
		.in_col (out_col_25_2),
		.out_row (out_row_26_2),
		.out_col (out_col_26_2),
		.out_data (out_data_26_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_3;
	wire signed [DATA_WIDTH-1:0] out_col_26_3;
	wire signed [DATA_WIDTH-1:0] out_data_26_3;
	integer_mac_pe mac_pe_26_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_2),
		.in_col (out_col_25_3),
		.out_row (out_row_26_3),
		.out_col (out_col_26_3),
		.out_data (out_data_26_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_4;
	wire signed [DATA_WIDTH-1:0] out_col_26_4;
	wire signed [DATA_WIDTH-1:0] out_data_26_4;
	integer_mac_pe mac_pe_26_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_3),
		.in_col (out_col_25_4),
		.out_row (out_row_26_4),
		.out_col (out_col_26_4),
		.out_data (out_data_26_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_5;
	wire signed [DATA_WIDTH-1:0] out_col_26_5;
	wire signed [DATA_WIDTH-1:0] out_data_26_5;
	integer_mac_pe mac_pe_26_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_4),
		.in_col (out_col_25_5),
		.out_row (out_row_26_5),
		.out_col (out_col_26_5),
		.out_data (out_data_26_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_6;
	wire signed [DATA_WIDTH-1:0] out_col_26_6;
	wire signed [DATA_WIDTH-1:0] out_data_26_6;
	integer_mac_pe mac_pe_26_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_5),
		.in_col (out_col_25_6),
		.out_row (out_row_26_6),
		.out_col (out_col_26_6),
		.out_data (out_data_26_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_7;
	wire signed [DATA_WIDTH-1:0] out_col_26_7;
	wire signed [DATA_WIDTH-1:0] out_data_26_7;
	integer_mac_pe mac_pe_26_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_6),
		.in_col (out_col_25_7),
		.out_row (out_row_26_7),
		.out_col (out_col_26_7),
		.out_data (out_data_26_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_8;
	wire signed [DATA_WIDTH-1:0] out_col_26_8;
	wire signed [DATA_WIDTH-1:0] out_data_26_8;
	integer_mac_pe mac_pe_26_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_7),
		.in_col (out_col_25_8),
		.out_row (out_row_26_8),
		.out_col (out_col_26_8),
		.out_data (out_data_26_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_9;
	wire signed [DATA_WIDTH-1:0] out_col_26_9;
	wire signed [DATA_WIDTH-1:0] out_data_26_9;
	integer_mac_pe mac_pe_26_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_8),
		.in_col (out_col_25_9),
		.out_row (out_row_26_9),
		.out_col (out_col_26_9),
		.out_data (out_data_26_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_10;
	wire signed [DATA_WIDTH-1:0] out_col_26_10;
	wire signed [DATA_WIDTH-1:0] out_data_26_10;
	integer_mac_pe mac_pe_26_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_9),
		.in_col (out_col_25_10),
		.out_row (out_row_26_10),
		.out_col (out_col_26_10),
		.out_data (out_data_26_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_11;
	wire signed [DATA_WIDTH-1:0] out_col_26_11;
	wire signed [DATA_WIDTH-1:0] out_data_26_11;
	integer_mac_pe mac_pe_26_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_10),
		.in_col (out_col_25_11),
		.out_row (out_row_26_11),
		.out_col (out_col_26_11),
		.out_data (out_data_26_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_12;
	wire signed [DATA_WIDTH-1:0] out_col_26_12;
	wire signed [DATA_WIDTH-1:0] out_data_26_12;
	integer_mac_pe mac_pe_26_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_11),
		.in_col (out_col_25_12),
		.out_row (out_row_26_12),
		.out_col (out_col_26_12),
		.out_data (out_data_26_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_13;
	wire signed [DATA_WIDTH-1:0] out_col_26_13;
	wire signed [DATA_WIDTH-1:0] out_data_26_13;
	integer_mac_pe mac_pe_26_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_12),
		.in_col (out_col_25_13),
		.out_row (out_row_26_13),
		.out_col (out_col_26_13),
		.out_data (out_data_26_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_14;
	wire signed [DATA_WIDTH-1:0] out_col_26_14;
	wire signed [DATA_WIDTH-1:0] out_data_26_14;
	integer_mac_pe mac_pe_26_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_13),
		.in_col (out_col_25_14),
		.out_row (out_row_26_14),
		.out_col (out_col_26_14),
		.out_data (out_data_26_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_15;
	wire signed [DATA_WIDTH-1:0] out_col_26_15;
	wire signed [DATA_WIDTH-1:0] out_data_26_15;
	integer_mac_pe mac_pe_26_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_14),
		.in_col (out_col_25_15),
		.out_row (out_row_26_15),
		.out_col (out_col_26_15),
		.out_data (out_data_26_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_16;
	wire signed [DATA_WIDTH-1:0] out_col_26_16;
	wire signed [DATA_WIDTH-1:0] out_data_26_16;
	integer_mac_pe mac_pe_26_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_15),
		.in_col (out_col_25_16),
		.out_row (out_row_26_16),
		.out_col (out_col_26_16),
		.out_data (out_data_26_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_17;
	wire signed [DATA_WIDTH-1:0] out_col_26_17;
	wire signed [DATA_WIDTH-1:0] out_data_26_17;
	integer_mac_pe mac_pe_26_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_16),
		.in_col (out_col_25_17),
		.out_row (out_row_26_17),
		.out_col (out_col_26_17),
		.out_data (out_data_26_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_18;
	wire signed [DATA_WIDTH-1:0] out_col_26_18;
	wire signed [DATA_WIDTH-1:0] out_data_26_18;
	integer_mac_pe mac_pe_26_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_17),
		.in_col (out_col_25_18),
		.out_row (out_row_26_18),
		.out_col (out_col_26_18),
		.out_data (out_data_26_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_19;
	wire signed [DATA_WIDTH-1:0] out_col_26_19;
	wire signed [DATA_WIDTH-1:0] out_data_26_19;
	integer_mac_pe mac_pe_26_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_18),
		.in_col (out_col_25_19),
		.out_row (out_row_26_19),
		.out_col (out_col_26_19),
		.out_data (out_data_26_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_20;
	wire signed [DATA_WIDTH-1:0] out_col_26_20;
	wire signed [DATA_WIDTH-1:0] out_data_26_20;
	integer_mac_pe mac_pe_26_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_19),
		.in_col (out_col_25_20),
		.out_row (out_row_26_20),
		.out_col (out_col_26_20),
		.out_data (out_data_26_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_21;
	wire signed [DATA_WIDTH-1:0] out_col_26_21;
	wire signed [DATA_WIDTH-1:0] out_data_26_21;
	integer_mac_pe mac_pe_26_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_20),
		.in_col (out_col_25_21),
		.out_row (out_row_26_21),
		.out_col (out_col_26_21),
		.out_data (out_data_26_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_22;
	wire signed [DATA_WIDTH-1:0] out_col_26_22;
	wire signed [DATA_WIDTH-1:0] out_data_26_22;
	integer_mac_pe mac_pe_26_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_21),
		.in_col (out_col_25_22),
		.out_row (out_row_26_22),
		.out_col (out_col_26_22),
		.out_data (out_data_26_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_23;
	wire signed [DATA_WIDTH-1:0] out_col_26_23;
	wire signed [DATA_WIDTH-1:0] out_data_26_23;
	integer_mac_pe mac_pe_26_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_22),
		.in_col (out_col_25_23),
		.out_row (out_row_26_23),
		.out_col (out_col_26_23),
		.out_data (out_data_26_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_24;
	wire signed [DATA_WIDTH-1:0] out_col_26_24;
	wire signed [DATA_WIDTH-1:0] out_data_26_24;
	integer_mac_pe mac_pe_26_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_23),
		.in_col (out_col_25_24),
		.out_row (out_row_26_24),
		.out_col (out_col_26_24),
		.out_data (out_data_26_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_25;
	wire signed [DATA_WIDTH-1:0] out_col_26_25;
	wire signed [DATA_WIDTH-1:0] out_data_26_25;
	integer_mac_pe mac_pe_26_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_24),
		.in_col (out_col_25_25),
		.out_row (out_row_26_25),
		.out_col (out_col_26_25),
		.out_data (out_data_26_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_26;
	wire signed [DATA_WIDTH-1:0] out_col_26_26;
	wire signed [DATA_WIDTH-1:0] out_data_26_26;
	integer_mac_pe mac_pe_26_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_25),
		.in_col (out_col_25_26),
		.out_row (out_row_26_26),
		.out_col (out_col_26_26),
		.out_data (out_data_26_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_27;
	wire signed [DATA_WIDTH-1:0] out_col_26_27;
	wire signed [DATA_WIDTH-1:0] out_data_26_27;
	integer_mac_pe mac_pe_26_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_26),
		.in_col (out_col_25_27),
		.out_row (out_row_26_27),
		.out_col (out_col_26_27),
		.out_data (out_data_26_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_28;
	wire signed [DATA_WIDTH-1:0] out_col_26_28;
	wire signed [DATA_WIDTH-1:0] out_data_26_28;
	integer_mac_pe mac_pe_26_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_27),
		.in_col (out_col_25_28),
		.out_row (out_row_26_28),
		.out_col (out_col_26_28),
		.out_data (out_data_26_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_29;
	wire signed [DATA_WIDTH-1:0] out_col_26_29;
	wire signed [DATA_WIDTH-1:0] out_data_26_29;
	integer_mac_pe mac_pe_26_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_28),
		.in_col (out_col_25_29),
		.out_row (out_row_26_29),
		.out_col (out_col_26_29),
		.out_data (out_data_26_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_30;
	wire signed [DATA_WIDTH-1:0] out_col_26_30;
	wire signed [DATA_WIDTH-1:0] out_data_26_30;
	integer_mac_pe mac_pe_26_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_29),
		.in_col (out_col_25_30),
		.out_row (out_row_26_30),
		.out_col (out_col_26_30),
		.out_data (out_data_26_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_26_31;
	wire signed [DATA_WIDTH-1:0] out_col_26_31;
	wire signed [DATA_WIDTH-1:0] out_data_26_31;
	integer_mac_pe mac_pe_26_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_26_30),
		.in_col (out_col_25_31),
		.out_row (out_row_26_31),
		.out_col (out_col_26_31),
		.out_data (out_data_26_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_0;
	wire signed [DATA_WIDTH-1:0] out_col_27_0;
	wire signed [DATA_WIDTH-1:0] out_data_27_0;
	integer_mac_pe mac_pe_27_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_27_out),
		.in_col (out_col_26_0),
		.out_row (out_row_27_0),
		.out_col (out_col_27_0),
		.out_data (out_data_27_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_1;
	wire signed [DATA_WIDTH-1:0] out_col_27_1;
	wire signed [DATA_WIDTH-1:0] out_data_27_1;
	integer_mac_pe mac_pe_27_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_0),
		.in_col (out_col_26_1),
		.out_row (out_row_27_1),
		.out_col (out_col_27_1),
		.out_data (out_data_27_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_2;
	wire signed [DATA_WIDTH-1:0] out_col_27_2;
	wire signed [DATA_WIDTH-1:0] out_data_27_2;
	integer_mac_pe mac_pe_27_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_1),
		.in_col (out_col_26_2),
		.out_row (out_row_27_2),
		.out_col (out_col_27_2),
		.out_data (out_data_27_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_3;
	wire signed [DATA_WIDTH-1:0] out_col_27_3;
	wire signed [DATA_WIDTH-1:0] out_data_27_3;
	integer_mac_pe mac_pe_27_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_2),
		.in_col (out_col_26_3),
		.out_row (out_row_27_3),
		.out_col (out_col_27_3),
		.out_data (out_data_27_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_4;
	wire signed [DATA_WIDTH-1:0] out_col_27_4;
	wire signed [DATA_WIDTH-1:0] out_data_27_4;
	integer_mac_pe mac_pe_27_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_3),
		.in_col (out_col_26_4),
		.out_row (out_row_27_4),
		.out_col (out_col_27_4),
		.out_data (out_data_27_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_5;
	wire signed [DATA_WIDTH-1:0] out_col_27_5;
	wire signed [DATA_WIDTH-1:0] out_data_27_5;
	integer_mac_pe mac_pe_27_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_4),
		.in_col (out_col_26_5),
		.out_row (out_row_27_5),
		.out_col (out_col_27_5),
		.out_data (out_data_27_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_6;
	wire signed [DATA_WIDTH-1:0] out_col_27_6;
	wire signed [DATA_WIDTH-1:0] out_data_27_6;
	integer_mac_pe mac_pe_27_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_5),
		.in_col (out_col_26_6),
		.out_row (out_row_27_6),
		.out_col (out_col_27_6),
		.out_data (out_data_27_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_7;
	wire signed [DATA_WIDTH-1:0] out_col_27_7;
	wire signed [DATA_WIDTH-1:0] out_data_27_7;
	integer_mac_pe mac_pe_27_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_6),
		.in_col (out_col_26_7),
		.out_row (out_row_27_7),
		.out_col (out_col_27_7),
		.out_data (out_data_27_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_8;
	wire signed [DATA_WIDTH-1:0] out_col_27_8;
	wire signed [DATA_WIDTH-1:0] out_data_27_8;
	integer_mac_pe mac_pe_27_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_7),
		.in_col (out_col_26_8),
		.out_row (out_row_27_8),
		.out_col (out_col_27_8),
		.out_data (out_data_27_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_9;
	wire signed [DATA_WIDTH-1:0] out_col_27_9;
	wire signed [DATA_WIDTH-1:0] out_data_27_9;
	integer_mac_pe mac_pe_27_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_8),
		.in_col (out_col_26_9),
		.out_row (out_row_27_9),
		.out_col (out_col_27_9),
		.out_data (out_data_27_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_10;
	wire signed [DATA_WIDTH-1:0] out_col_27_10;
	wire signed [DATA_WIDTH-1:0] out_data_27_10;
	integer_mac_pe mac_pe_27_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_9),
		.in_col (out_col_26_10),
		.out_row (out_row_27_10),
		.out_col (out_col_27_10),
		.out_data (out_data_27_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_11;
	wire signed [DATA_WIDTH-1:0] out_col_27_11;
	wire signed [DATA_WIDTH-1:0] out_data_27_11;
	integer_mac_pe mac_pe_27_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_10),
		.in_col (out_col_26_11),
		.out_row (out_row_27_11),
		.out_col (out_col_27_11),
		.out_data (out_data_27_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_12;
	wire signed [DATA_WIDTH-1:0] out_col_27_12;
	wire signed [DATA_WIDTH-1:0] out_data_27_12;
	integer_mac_pe mac_pe_27_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_11),
		.in_col (out_col_26_12),
		.out_row (out_row_27_12),
		.out_col (out_col_27_12),
		.out_data (out_data_27_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_13;
	wire signed [DATA_WIDTH-1:0] out_col_27_13;
	wire signed [DATA_WIDTH-1:0] out_data_27_13;
	integer_mac_pe mac_pe_27_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_12),
		.in_col (out_col_26_13),
		.out_row (out_row_27_13),
		.out_col (out_col_27_13),
		.out_data (out_data_27_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_14;
	wire signed [DATA_WIDTH-1:0] out_col_27_14;
	wire signed [DATA_WIDTH-1:0] out_data_27_14;
	integer_mac_pe mac_pe_27_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_13),
		.in_col (out_col_26_14),
		.out_row (out_row_27_14),
		.out_col (out_col_27_14),
		.out_data (out_data_27_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_15;
	wire signed [DATA_WIDTH-1:0] out_col_27_15;
	wire signed [DATA_WIDTH-1:0] out_data_27_15;
	integer_mac_pe mac_pe_27_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_14),
		.in_col (out_col_26_15),
		.out_row (out_row_27_15),
		.out_col (out_col_27_15),
		.out_data (out_data_27_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_16;
	wire signed [DATA_WIDTH-1:0] out_col_27_16;
	wire signed [DATA_WIDTH-1:0] out_data_27_16;
	integer_mac_pe mac_pe_27_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_15),
		.in_col (out_col_26_16),
		.out_row (out_row_27_16),
		.out_col (out_col_27_16),
		.out_data (out_data_27_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_17;
	wire signed [DATA_WIDTH-1:0] out_col_27_17;
	wire signed [DATA_WIDTH-1:0] out_data_27_17;
	integer_mac_pe mac_pe_27_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_16),
		.in_col (out_col_26_17),
		.out_row (out_row_27_17),
		.out_col (out_col_27_17),
		.out_data (out_data_27_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_18;
	wire signed [DATA_WIDTH-1:0] out_col_27_18;
	wire signed [DATA_WIDTH-1:0] out_data_27_18;
	integer_mac_pe mac_pe_27_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_17),
		.in_col (out_col_26_18),
		.out_row (out_row_27_18),
		.out_col (out_col_27_18),
		.out_data (out_data_27_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_19;
	wire signed [DATA_WIDTH-1:0] out_col_27_19;
	wire signed [DATA_WIDTH-1:0] out_data_27_19;
	integer_mac_pe mac_pe_27_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_18),
		.in_col (out_col_26_19),
		.out_row (out_row_27_19),
		.out_col (out_col_27_19),
		.out_data (out_data_27_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_20;
	wire signed [DATA_WIDTH-1:0] out_col_27_20;
	wire signed [DATA_WIDTH-1:0] out_data_27_20;
	integer_mac_pe mac_pe_27_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_19),
		.in_col (out_col_26_20),
		.out_row (out_row_27_20),
		.out_col (out_col_27_20),
		.out_data (out_data_27_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_21;
	wire signed [DATA_WIDTH-1:0] out_col_27_21;
	wire signed [DATA_WIDTH-1:0] out_data_27_21;
	integer_mac_pe mac_pe_27_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_20),
		.in_col (out_col_26_21),
		.out_row (out_row_27_21),
		.out_col (out_col_27_21),
		.out_data (out_data_27_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_22;
	wire signed [DATA_WIDTH-1:0] out_col_27_22;
	wire signed [DATA_WIDTH-1:0] out_data_27_22;
	integer_mac_pe mac_pe_27_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_21),
		.in_col (out_col_26_22),
		.out_row (out_row_27_22),
		.out_col (out_col_27_22),
		.out_data (out_data_27_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_23;
	wire signed [DATA_WIDTH-1:0] out_col_27_23;
	wire signed [DATA_WIDTH-1:0] out_data_27_23;
	integer_mac_pe mac_pe_27_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_22),
		.in_col (out_col_26_23),
		.out_row (out_row_27_23),
		.out_col (out_col_27_23),
		.out_data (out_data_27_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_24;
	wire signed [DATA_WIDTH-1:0] out_col_27_24;
	wire signed [DATA_WIDTH-1:0] out_data_27_24;
	integer_mac_pe mac_pe_27_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_23),
		.in_col (out_col_26_24),
		.out_row (out_row_27_24),
		.out_col (out_col_27_24),
		.out_data (out_data_27_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_25;
	wire signed [DATA_WIDTH-1:0] out_col_27_25;
	wire signed [DATA_WIDTH-1:0] out_data_27_25;
	integer_mac_pe mac_pe_27_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_24),
		.in_col (out_col_26_25),
		.out_row (out_row_27_25),
		.out_col (out_col_27_25),
		.out_data (out_data_27_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_26;
	wire signed [DATA_WIDTH-1:0] out_col_27_26;
	wire signed [DATA_WIDTH-1:0] out_data_27_26;
	integer_mac_pe mac_pe_27_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_25),
		.in_col (out_col_26_26),
		.out_row (out_row_27_26),
		.out_col (out_col_27_26),
		.out_data (out_data_27_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_27;
	wire signed [DATA_WIDTH-1:0] out_col_27_27;
	wire signed [DATA_WIDTH-1:0] out_data_27_27;
	integer_mac_pe mac_pe_27_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_26),
		.in_col (out_col_26_27),
		.out_row (out_row_27_27),
		.out_col (out_col_27_27),
		.out_data (out_data_27_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_28;
	wire signed [DATA_WIDTH-1:0] out_col_27_28;
	wire signed [DATA_WIDTH-1:0] out_data_27_28;
	integer_mac_pe mac_pe_27_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_27),
		.in_col (out_col_26_28),
		.out_row (out_row_27_28),
		.out_col (out_col_27_28),
		.out_data (out_data_27_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_29;
	wire signed [DATA_WIDTH-1:0] out_col_27_29;
	wire signed [DATA_WIDTH-1:0] out_data_27_29;
	integer_mac_pe mac_pe_27_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_28),
		.in_col (out_col_26_29),
		.out_row (out_row_27_29),
		.out_col (out_col_27_29),
		.out_data (out_data_27_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_30;
	wire signed [DATA_WIDTH-1:0] out_col_27_30;
	wire signed [DATA_WIDTH-1:0] out_data_27_30;
	integer_mac_pe mac_pe_27_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_29),
		.in_col (out_col_26_30),
		.out_row (out_row_27_30),
		.out_col (out_col_27_30),
		.out_data (out_data_27_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_27_31;
	wire signed [DATA_WIDTH-1:0] out_col_27_31;
	wire signed [DATA_WIDTH-1:0] out_data_27_31;
	integer_mac_pe mac_pe_27_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_27_30),
		.in_col (out_col_26_31),
		.out_row (out_row_27_31),
		.out_col (out_col_27_31),
		.out_data (out_data_27_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_0;
	wire signed [DATA_WIDTH-1:0] out_col_28_0;
	wire signed [DATA_WIDTH-1:0] out_data_28_0;
	integer_mac_pe mac_pe_28_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_28_out),
		.in_col (out_col_27_0),
		.out_row (out_row_28_0),
		.out_col (out_col_28_0),
		.out_data (out_data_28_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_1;
	wire signed [DATA_WIDTH-1:0] out_col_28_1;
	wire signed [DATA_WIDTH-1:0] out_data_28_1;
	integer_mac_pe mac_pe_28_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_0),
		.in_col (out_col_27_1),
		.out_row (out_row_28_1),
		.out_col (out_col_28_1),
		.out_data (out_data_28_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_2;
	wire signed [DATA_WIDTH-1:0] out_col_28_2;
	wire signed [DATA_WIDTH-1:0] out_data_28_2;
	integer_mac_pe mac_pe_28_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_1),
		.in_col (out_col_27_2),
		.out_row (out_row_28_2),
		.out_col (out_col_28_2),
		.out_data (out_data_28_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_3;
	wire signed [DATA_WIDTH-1:0] out_col_28_3;
	wire signed [DATA_WIDTH-1:0] out_data_28_3;
	integer_mac_pe mac_pe_28_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_2),
		.in_col (out_col_27_3),
		.out_row (out_row_28_3),
		.out_col (out_col_28_3),
		.out_data (out_data_28_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_4;
	wire signed [DATA_WIDTH-1:0] out_col_28_4;
	wire signed [DATA_WIDTH-1:0] out_data_28_4;
	integer_mac_pe mac_pe_28_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_3),
		.in_col (out_col_27_4),
		.out_row (out_row_28_4),
		.out_col (out_col_28_4),
		.out_data (out_data_28_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_5;
	wire signed [DATA_WIDTH-1:0] out_col_28_5;
	wire signed [DATA_WIDTH-1:0] out_data_28_5;
	integer_mac_pe mac_pe_28_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_4),
		.in_col (out_col_27_5),
		.out_row (out_row_28_5),
		.out_col (out_col_28_5),
		.out_data (out_data_28_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_6;
	wire signed [DATA_WIDTH-1:0] out_col_28_6;
	wire signed [DATA_WIDTH-1:0] out_data_28_6;
	integer_mac_pe mac_pe_28_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_5),
		.in_col (out_col_27_6),
		.out_row (out_row_28_6),
		.out_col (out_col_28_6),
		.out_data (out_data_28_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_7;
	wire signed [DATA_WIDTH-1:0] out_col_28_7;
	wire signed [DATA_WIDTH-1:0] out_data_28_7;
	integer_mac_pe mac_pe_28_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_6),
		.in_col (out_col_27_7),
		.out_row (out_row_28_7),
		.out_col (out_col_28_7),
		.out_data (out_data_28_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_8;
	wire signed [DATA_WIDTH-1:0] out_col_28_8;
	wire signed [DATA_WIDTH-1:0] out_data_28_8;
	integer_mac_pe mac_pe_28_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_7),
		.in_col (out_col_27_8),
		.out_row (out_row_28_8),
		.out_col (out_col_28_8),
		.out_data (out_data_28_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_9;
	wire signed [DATA_WIDTH-1:0] out_col_28_9;
	wire signed [DATA_WIDTH-1:0] out_data_28_9;
	integer_mac_pe mac_pe_28_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_8),
		.in_col (out_col_27_9),
		.out_row (out_row_28_9),
		.out_col (out_col_28_9),
		.out_data (out_data_28_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_10;
	wire signed [DATA_WIDTH-1:0] out_col_28_10;
	wire signed [DATA_WIDTH-1:0] out_data_28_10;
	integer_mac_pe mac_pe_28_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_9),
		.in_col (out_col_27_10),
		.out_row (out_row_28_10),
		.out_col (out_col_28_10),
		.out_data (out_data_28_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_11;
	wire signed [DATA_WIDTH-1:0] out_col_28_11;
	wire signed [DATA_WIDTH-1:0] out_data_28_11;
	integer_mac_pe mac_pe_28_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_10),
		.in_col (out_col_27_11),
		.out_row (out_row_28_11),
		.out_col (out_col_28_11),
		.out_data (out_data_28_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_12;
	wire signed [DATA_WIDTH-1:0] out_col_28_12;
	wire signed [DATA_WIDTH-1:0] out_data_28_12;
	integer_mac_pe mac_pe_28_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_11),
		.in_col (out_col_27_12),
		.out_row (out_row_28_12),
		.out_col (out_col_28_12),
		.out_data (out_data_28_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_13;
	wire signed [DATA_WIDTH-1:0] out_col_28_13;
	wire signed [DATA_WIDTH-1:0] out_data_28_13;
	integer_mac_pe mac_pe_28_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_12),
		.in_col (out_col_27_13),
		.out_row (out_row_28_13),
		.out_col (out_col_28_13),
		.out_data (out_data_28_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_14;
	wire signed [DATA_WIDTH-1:0] out_col_28_14;
	wire signed [DATA_WIDTH-1:0] out_data_28_14;
	integer_mac_pe mac_pe_28_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_13),
		.in_col (out_col_27_14),
		.out_row (out_row_28_14),
		.out_col (out_col_28_14),
		.out_data (out_data_28_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_15;
	wire signed [DATA_WIDTH-1:0] out_col_28_15;
	wire signed [DATA_WIDTH-1:0] out_data_28_15;
	integer_mac_pe mac_pe_28_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_14),
		.in_col (out_col_27_15),
		.out_row (out_row_28_15),
		.out_col (out_col_28_15),
		.out_data (out_data_28_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_16;
	wire signed [DATA_WIDTH-1:0] out_col_28_16;
	wire signed [DATA_WIDTH-1:0] out_data_28_16;
	integer_mac_pe mac_pe_28_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_15),
		.in_col (out_col_27_16),
		.out_row (out_row_28_16),
		.out_col (out_col_28_16),
		.out_data (out_data_28_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_17;
	wire signed [DATA_WIDTH-1:0] out_col_28_17;
	wire signed [DATA_WIDTH-1:0] out_data_28_17;
	integer_mac_pe mac_pe_28_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_16),
		.in_col (out_col_27_17),
		.out_row (out_row_28_17),
		.out_col (out_col_28_17),
		.out_data (out_data_28_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_18;
	wire signed [DATA_WIDTH-1:0] out_col_28_18;
	wire signed [DATA_WIDTH-1:0] out_data_28_18;
	integer_mac_pe mac_pe_28_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_17),
		.in_col (out_col_27_18),
		.out_row (out_row_28_18),
		.out_col (out_col_28_18),
		.out_data (out_data_28_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_19;
	wire signed [DATA_WIDTH-1:0] out_col_28_19;
	wire signed [DATA_WIDTH-1:0] out_data_28_19;
	integer_mac_pe mac_pe_28_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_18),
		.in_col (out_col_27_19),
		.out_row (out_row_28_19),
		.out_col (out_col_28_19),
		.out_data (out_data_28_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_20;
	wire signed [DATA_WIDTH-1:0] out_col_28_20;
	wire signed [DATA_WIDTH-1:0] out_data_28_20;
	integer_mac_pe mac_pe_28_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_19),
		.in_col (out_col_27_20),
		.out_row (out_row_28_20),
		.out_col (out_col_28_20),
		.out_data (out_data_28_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_21;
	wire signed [DATA_WIDTH-1:0] out_col_28_21;
	wire signed [DATA_WIDTH-1:0] out_data_28_21;
	integer_mac_pe mac_pe_28_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_20),
		.in_col (out_col_27_21),
		.out_row (out_row_28_21),
		.out_col (out_col_28_21),
		.out_data (out_data_28_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_22;
	wire signed [DATA_WIDTH-1:0] out_col_28_22;
	wire signed [DATA_WIDTH-1:0] out_data_28_22;
	integer_mac_pe mac_pe_28_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_21),
		.in_col (out_col_27_22),
		.out_row (out_row_28_22),
		.out_col (out_col_28_22),
		.out_data (out_data_28_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_23;
	wire signed [DATA_WIDTH-1:0] out_col_28_23;
	wire signed [DATA_WIDTH-1:0] out_data_28_23;
	integer_mac_pe mac_pe_28_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_22),
		.in_col (out_col_27_23),
		.out_row (out_row_28_23),
		.out_col (out_col_28_23),
		.out_data (out_data_28_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_24;
	wire signed [DATA_WIDTH-1:0] out_col_28_24;
	wire signed [DATA_WIDTH-1:0] out_data_28_24;
	integer_mac_pe mac_pe_28_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_23),
		.in_col (out_col_27_24),
		.out_row (out_row_28_24),
		.out_col (out_col_28_24),
		.out_data (out_data_28_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_25;
	wire signed [DATA_WIDTH-1:0] out_col_28_25;
	wire signed [DATA_WIDTH-1:0] out_data_28_25;
	integer_mac_pe mac_pe_28_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_24),
		.in_col (out_col_27_25),
		.out_row (out_row_28_25),
		.out_col (out_col_28_25),
		.out_data (out_data_28_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_26;
	wire signed [DATA_WIDTH-1:0] out_col_28_26;
	wire signed [DATA_WIDTH-1:0] out_data_28_26;
	integer_mac_pe mac_pe_28_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_25),
		.in_col (out_col_27_26),
		.out_row (out_row_28_26),
		.out_col (out_col_28_26),
		.out_data (out_data_28_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_27;
	wire signed [DATA_WIDTH-1:0] out_col_28_27;
	wire signed [DATA_WIDTH-1:0] out_data_28_27;
	integer_mac_pe mac_pe_28_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_26),
		.in_col (out_col_27_27),
		.out_row (out_row_28_27),
		.out_col (out_col_28_27),
		.out_data (out_data_28_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_28;
	wire signed [DATA_WIDTH-1:0] out_col_28_28;
	wire signed [DATA_WIDTH-1:0] out_data_28_28;
	integer_mac_pe mac_pe_28_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_27),
		.in_col (out_col_27_28),
		.out_row (out_row_28_28),
		.out_col (out_col_28_28),
		.out_data (out_data_28_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_29;
	wire signed [DATA_WIDTH-1:0] out_col_28_29;
	wire signed [DATA_WIDTH-1:0] out_data_28_29;
	integer_mac_pe mac_pe_28_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_28),
		.in_col (out_col_27_29),
		.out_row (out_row_28_29),
		.out_col (out_col_28_29),
		.out_data (out_data_28_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_30;
	wire signed [DATA_WIDTH-1:0] out_col_28_30;
	wire signed [DATA_WIDTH-1:0] out_data_28_30;
	integer_mac_pe mac_pe_28_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_29),
		.in_col (out_col_27_30),
		.out_row (out_row_28_30),
		.out_col (out_col_28_30),
		.out_data (out_data_28_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_28_31;
	wire signed [DATA_WIDTH-1:0] out_col_28_31;
	wire signed [DATA_WIDTH-1:0] out_data_28_31;
	integer_mac_pe mac_pe_28_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_28_30),
		.in_col (out_col_27_31),
		.out_row (out_row_28_31),
		.out_col (out_col_28_31),
		.out_data (out_data_28_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_0;
	wire signed [DATA_WIDTH-1:0] out_col_29_0;
	wire signed [DATA_WIDTH-1:0] out_data_29_0;
	integer_mac_pe mac_pe_29_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_29_out),
		.in_col (out_col_28_0),
		.out_row (out_row_29_0),
		.out_col (out_col_29_0),
		.out_data (out_data_29_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_1;
	wire signed [DATA_WIDTH-1:0] out_col_29_1;
	wire signed [DATA_WIDTH-1:0] out_data_29_1;
	integer_mac_pe mac_pe_29_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_0),
		.in_col (out_col_28_1),
		.out_row (out_row_29_1),
		.out_col (out_col_29_1),
		.out_data (out_data_29_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_2;
	wire signed [DATA_WIDTH-1:0] out_col_29_2;
	wire signed [DATA_WIDTH-1:0] out_data_29_2;
	integer_mac_pe mac_pe_29_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_1),
		.in_col (out_col_28_2),
		.out_row (out_row_29_2),
		.out_col (out_col_29_2),
		.out_data (out_data_29_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_3;
	wire signed [DATA_WIDTH-1:0] out_col_29_3;
	wire signed [DATA_WIDTH-1:0] out_data_29_3;
	integer_mac_pe mac_pe_29_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_2),
		.in_col (out_col_28_3),
		.out_row (out_row_29_3),
		.out_col (out_col_29_3),
		.out_data (out_data_29_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_4;
	wire signed [DATA_WIDTH-1:0] out_col_29_4;
	wire signed [DATA_WIDTH-1:0] out_data_29_4;
	integer_mac_pe mac_pe_29_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_3),
		.in_col (out_col_28_4),
		.out_row (out_row_29_4),
		.out_col (out_col_29_4),
		.out_data (out_data_29_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_5;
	wire signed [DATA_WIDTH-1:0] out_col_29_5;
	wire signed [DATA_WIDTH-1:0] out_data_29_5;
	integer_mac_pe mac_pe_29_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_4),
		.in_col (out_col_28_5),
		.out_row (out_row_29_5),
		.out_col (out_col_29_5),
		.out_data (out_data_29_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_6;
	wire signed [DATA_WIDTH-1:0] out_col_29_6;
	wire signed [DATA_WIDTH-1:0] out_data_29_6;
	integer_mac_pe mac_pe_29_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_5),
		.in_col (out_col_28_6),
		.out_row (out_row_29_6),
		.out_col (out_col_29_6),
		.out_data (out_data_29_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_7;
	wire signed [DATA_WIDTH-1:0] out_col_29_7;
	wire signed [DATA_WIDTH-1:0] out_data_29_7;
	integer_mac_pe mac_pe_29_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_6),
		.in_col (out_col_28_7),
		.out_row (out_row_29_7),
		.out_col (out_col_29_7),
		.out_data (out_data_29_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_8;
	wire signed [DATA_WIDTH-1:0] out_col_29_8;
	wire signed [DATA_WIDTH-1:0] out_data_29_8;
	integer_mac_pe mac_pe_29_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_7),
		.in_col (out_col_28_8),
		.out_row (out_row_29_8),
		.out_col (out_col_29_8),
		.out_data (out_data_29_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_9;
	wire signed [DATA_WIDTH-1:0] out_col_29_9;
	wire signed [DATA_WIDTH-1:0] out_data_29_9;
	integer_mac_pe mac_pe_29_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_8),
		.in_col (out_col_28_9),
		.out_row (out_row_29_9),
		.out_col (out_col_29_9),
		.out_data (out_data_29_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_10;
	wire signed [DATA_WIDTH-1:0] out_col_29_10;
	wire signed [DATA_WIDTH-1:0] out_data_29_10;
	integer_mac_pe mac_pe_29_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_9),
		.in_col (out_col_28_10),
		.out_row (out_row_29_10),
		.out_col (out_col_29_10),
		.out_data (out_data_29_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_11;
	wire signed [DATA_WIDTH-1:0] out_col_29_11;
	wire signed [DATA_WIDTH-1:0] out_data_29_11;
	integer_mac_pe mac_pe_29_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_10),
		.in_col (out_col_28_11),
		.out_row (out_row_29_11),
		.out_col (out_col_29_11),
		.out_data (out_data_29_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_12;
	wire signed [DATA_WIDTH-1:0] out_col_29_12;
	wire signed [DATA_WIDTH-1:0] out_data_29_12;
	integer_mac_pe mac_pe_29_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_11),
		.in_col (out_col_28_12),
		.out_row (out_row_29_12),
		.out_col (out_col_29_12),
		.out_data (out_data_29_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_13;
	wire signed [DATA_WIDTH-1:0] out_col_29_13;
	wire signed [DATA_WIDTH-1:0] out_data_29_13;
	integer_mac_pe mac_pe_29_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_12),
		.in_col (out_col_28_13),
		.out_row (out_row_29_13),
		.out_col (out_col_29_13),
		.out_data (out_data_29_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_14;
	wire signed [DATA_WIDTH-1:0] out_col_29_14;
	wire signed [DATA_WIDTH-1:0] out_data_29_14;
	integer_mac_pe mac_pe_29_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_13),
		.in_col (out_col_28_14),
		.out_row (out_row_29_14),
		.out_col (out_col_29_14),
		.out_data (out_data_29_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_15;
	wire signed [DATA_WIDTH-1:0] out_col_29_15;
	wire signed [DATA_WIDTH-1:0] out_data_29_15;
	integer_mac_pe mac_pe_29_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_14),
		.in_col (out_col_28_15),
		.out_row (out_row_29_15),
		.out_col (out_col_29_15),
		.out_data (out_data_29_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_16;
	wire signed [DATA_WIDTH-1:0] out_col_29_16;
	wire signed [DATA_WIDTH-1:0] out_data_29_16;
	integer_mac_pe mac_pe_29_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_15),
		.in_col (out_col_28_16),
		.out_row (out_row_29_16),
		.out_col (out_col_29_16),
		.out_data (out_data_29_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_17;
	wire signed [DATA_WIDTH-1:0] out_col_29_17;
	wire signed [DATA_WIDTH-1:0] out_data_29_17;
	integer_mac_pe mac_pe_29_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_16),
		.in_col (out_col_28_17),
		.out_row (out_row_29_17),
		.out_col (out_col_29_17),
		.out_data (out_data_29_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_18;
	wire signed [DATA_WIDTH-1:0] out_col_29_18;
	wire signed [DATA_WIDTH-1:0] out_data_29_18;
	integer_mac_pe mac_pe_29_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_17),
		.in_col (out_col_28_18),
		.out_row (out_row_29_18),
		.out_col (out_col_29_18),
		.out_data (out_data_29_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_19;
	wire signed [DATA_WIDTH-1:0] out_col_29_19;
	wire signed [DATA_WIDTH-1:0] out_data_29_19;
	integer_mac_pe mac_pe_29_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_18),
		.in_col (out_col_28_19),
		.out_row (out_row_29_19),
		.out_col (out_col_29_19),
		.out_data (out_data_29_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_20;
	wire signed [DATA_WIDTH-1:0] out_col_29_20;
	wire signed [DATA_WIDTH-1:0] out_data_29_20;
	integer_mac_pe mac_pe_29_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_19),
		.in_col (out_col_28_20),
		.out_row (out_row_29_20),
		.out_col (out_col_29_20),
		.out_data (out_data_29_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_21;
	wire signed [DATA_WIDTH-1:0] out_col_29_21;
	wire signed [DATA_WIDTH-1:0] out_data_29_21;
	integer_mac_pe mac_pe_29_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_20),
		.in_col (out_col_28_21),
		.out_row (out_row_29_21),
		.out_col (out_col_29_21),
		.out_data (out_data_29_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_22;
	wire signed [DATA_WIDTH-1:0] out_col_29_22;
	wire signed [DATA_WIDTH-1:0] out_data_29_22;
	integer_mac_pe mac_pe_29_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_21),
		.in_col (out_col_28_22),
		.out_row (out_row_29_22),
		.out_col (out_col_29_22),
		.out_data (out_data_29_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_23;
	wire signed [DATA_WIDTH-1:0] out_col_29_23;
	wire signed [DATA_WIDTH-1:0] out_data_29_23;
	integer_mac_pe mac_pe_29_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_22),
		.in_col (out_col_28_23),
		.out_row (out_row_29_23),
		.out_col (out_col_29_23),
		.out_data (out_data_29_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_24;
	wire signed [DATA_WIDTH-1:0] out_col_29_24;
	wire signed [DATA_WIDTH-1:0] out_data_29_24;
	integer_mac_pe mac_pe_29_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_23),
		.in_col (out_col_28_24),
		.out_row (out_row_29_24),
		.out_col (out_col_29_24),
		.out_data (out_data_29_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_25;
	wire signed [DATA_WIDTH-1:0] out_col_29_25;
	wire signed [DATA_WIDTH-1:0] out_data_29_25;
	integer_mac_pe mac_pe_29_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_24),
		.in_col (out_col_28_25),
		.out_row (out_row_29_25),
		.out_col (out_col_29_25),
		.out_data (out_data_29_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_26;
	wire signed [DATA_WIDTH-1:0] out_col_29_26;
	wire signed [DATA_WIDTH-1:0] out_data_29_26;
	integer_mac_pe mac_pe_29_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_25),
		.in_col (out_col_28_26),
		.out_row (out_row_29_26),
		.out_col (out_col_29_26),
		.out_data (out_data_29_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_27;
	wire signed [DATA_WIDTH-1:0] out_col_29_27;
	wire signed [DATA_WIDTH-1:0] out_data_29_27;
	integer_mac_pe mac_pe_29_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_26),
		.in_col (out_col_28_27),
		.out_row (out_row_29_27),
		.out_col (out_col_29_27),
		.out_data (out_data_29_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_28;
	wire signed [DATA_WIDTH-1:0] out_col_29_28;
	wire signed [DATA_WIDTH-1:0] out_data_29_28;
	integer_mac_pe mac_pe_29_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_27),
		.in_col (out_col_28_28),
		.out_row (out_row_29_28),
		.out_col (out_col_29_28),
		.out_data (out_data_29_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_29;
	wire signed [DATA_WIDTH-1:0] out_col_29_29;
	wire signed [DATA_WIDTH-1:0] out_data_29_29;
	integer_mac_pe mac_pe_29_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_28),
		.in_col (out_col_28_29),
		.out_row (out_row_29_29),
		.out_col (out_col_29_29),
		.out_data (out_data_29_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_30;
	wire signed [DATA_WIDTH-1:0] out_col_29_30;
	wire signed [DATA_WIDTH-1:0] out_data_29_30;
	integer_mac_pe mac_pe_29_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_29),
		.in_col (out_col_28_30),
		.out_row (out_row_29_30),
		.out_col (out_col_29_30),
		.out_data (out_data_29_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_29_31;
	wire signed [DATA_WIDTH-1:0] out_col_29_31;
	wire signed [DATA_WIDTH-1:0] out_data_29_31;
	integer_mac_pe mac_pe_29_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_29_30),
		.in_col (out_col_28_31),
		.out_row (out_row_29_31),
		.out_col (out_col_29_31),
		.out_data (out_data_29_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_0;
	wire signed [DATA_WIDTH-1:0] out_col_30_0;
	wire signed [DATA_WIDTH-1:0] out_data_30_0;
	integer_mac_pe mac_pe_30_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_30_out),
		.in_col (out_col_29_0),
		.out_row (out_row_30_0),
		.out_col (out_col_30_0),
		.out_data (out_data_30_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_1;
	wire signed [DATA_WIDTH-1:0] out_col_30_1;
	wire signed [DATA_WIDTH-1:0] out_data_30_1;
	integer_mac_pe mac_pe_30_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_0),
		.in_col (out_col_29_1),
		.out_row (out_row_30_1),
		.out_col (out_col_30_1),
		.out_data (out_data_30_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_2;
	wire signed [DATA_WIDTH-1:0] out_col_30_2;
	wire signed [DATA_WIDTH-1:0] out_data_30_2;
	integer_mac_pe mac_pe_30_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_1),
		.in_col (out_col_29_2),
		.out_row (out_row_30_2),
		.out_col (out_col_30_2),
		.out_data (out_data_30_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_3;
	wire signed [DATA_WIDTH-1:0] out_col_30_3;
	wire signed [DATA_WIDTH-1:0] out_data_30_3;
	integer_mac_pe mac_pe_30_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_2),
		.in_col (out_col_29_3),
		.out_row (out_row_30_3),
		.out_col (out_col_30_3),
		.out_data (out_data_30_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_4;
	wire signed [DATA_WIDTH-1:0] out_col_30_4;
	wire signed [DATA_WIDTH-1:0] out_data_30_4;
	integer_mac_pe mac_pe_30_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_3),
		.in_col (out_col_29_4),
		.out_row (out_row_30_4),
		.out_col (out_col_30_4),
		.out_data (out_data_30_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_5;
	wire signed [DATA_WIDTH-1:0] out_col_30_5;
	wire signed [DATA_WIDTH-1:0] out_data_30_5;
	integer_mac_pe mac_pe_30_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_4),
		.in_col (out_col_29_5),
		.out_row (out_row_30_5),
		.out_col (out_col_30_5),
		.out_data (out_data_30_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_6;
	wire signed [DATA_WIDTH-1:0] out_col_30_6;
	wire signed [DATA_WIDTH-1:0] out_data_30_6;
	integer_mac_pe mac_pe_30_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_5),
		.in_col (out_col_29_6),
		.out_row (out_row_30_6),
		.out_col (out_col_30_6),
		.out_data (out_data_30_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_7;
	wire signed [DATA_WIDTH-1:0] out_col_30_7;
	wire signed [DATA_WIDTH-1:0] out_data_30_7;
	integer_mac_pe mac_pe_30_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_6),
		.in_col (out_col_29_7),
		.out_row (out_row_30_7),
		.out_col (out_col_30_7),
		.out_data (out_data_30_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_8;
	wire signed [DATA_WIDTH-1:0] out_col_30_8;
	wire signed [DATA_WIDTH-1:0] out_data_30_8;
	integer_mac_pe mac_pe_30_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_7),
		.in_col (out_col_29_8),
		.out_row (out_row_30_8),
		.out_col (out_col_30_8),
		.out_data (out_data_30_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_9;
	wire signed [DATA_WIDTH-1:0] out_col_30_9;
	wire signed [DATA_WIDTH-1:0] out_data_30_9;
	integer_mac_pe mac_pe_30_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_8),
		.in_col (out_col_29_9),
		.out_row (out_row_30_9),
		.out_col (out_col_30_9),
		.out_data (out_data_30_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_10;
	wire signed [DATA_WIDTH-1:0] out_col_30_10;
	wire signed [DATA_WIDTH-1:0] out_data_30_10;
	integer_mac_pe mac_pe_30_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_9),
		.in_col (out_col_29_10),
		.out_row (out_row_30_10),
		.out_col (out_col_30_10),
		.out_data (out_data_30_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_11;
	wire signed [DATA_WIDTH-1:0] out_col_30_11;
	wire signed [DATA_WIDTH-1:0] out_data_30_11;
	integer_mac_pe mac_pe_30_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_10),
		.in_col (out_col_29_11),
		.out_row (out_row_30_11),
		.out_col (out_col_30_11),
		.out_data (out_data_30_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_12;
	wire signed [DATA_WIDTH-1:0] out_col_30_12;
	wire signed [DATA_WIDTH-1:0] out_data_30_12;
	integer_mac_pe mac_pe_30_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_11),
		.in_col (out_col_29_12),
		.out_row (out_row_30_12),
		.out_col (out_col_30_12),
		.out_data (out_data_30_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_13;
	wire signed [DATA_WIDTH-1:0] out_col_30_13;
	wire signed [DATA_WIDTH-1:0] out_data_30_13;
	integer_mac_pe mac_pe_30_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_12),
		.in_col (out_col_29_13),
		.out_row (out_row_30_13),
		.out_col (out_col_30_13),
		.out_data (out_data_30_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_14;
	wire signed [DATA_WIDTH-1:0] out_col_30_14;
	wire signed [DATA_WIDTH-1:0] out_data_30_14;
	integer_mac_pe mac_pe_30_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_13),
		.in_col (out_col_29_14),
		.out_row (out_row_30_14),
		.out_col (out_col_30_14),
		.out_data (out_data_30_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_15;
	wire signed [DATA_WIDTH-1:0] out_col_30_15;
	wire signed [DATA_WIDTH-1:0] out_data_30_15;
	integer_mac_pe mac_pe_30_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_14),
		.in_col (out_col_29_15),
		.out_row (out_row_30_15),
		.out_col (out_col_30_15),
		.out_data (out_data_30_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_16;
	wire signed [DATA_WIDTH-1:0] out_col_30_16;
	wire signed [DATA_WIDTH-1:0] out_data_30_16;
	integer_mac_pe mac_pe_30_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_15),
		.in_col (out_col_29_16),
		.out_row (out_row_30_16),
		.out_col (out_col_30_16),
		.out_data (out_data_30_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_17;
	wire signed [DATA_WIDTH-1:0] out_col_30_17;
	wire signed [DATA_WIDTH-1:0] out_data_30_17;
	integer_mac_pe mac_pe_30_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_16),
		.in_col (out_col_29_17),
		.out_row (out_row_30_17),
		.out_col (out_col_30_17),
		.out_data (out_data_30_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_18;
	wire signed [DATA_WIDTH-1:0] out_col_30_18;
	wire signed [DATA_WIDTH-1:0] out_data_30_18;
	integer_mac_pe mac_pe_30_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_17),
		.in_col (out_col_29_18),
		.out_row (out_row_30_18),
		.out_col (out_col_30_18),
		.out_data (out_data_30_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_19;
	wire signed [DATA_WIDTH-1:0] out_col_30_19;
	wire signed [DATA_WIDTH-1:0] out_data_30_19;
	integer_mac_pe mac_pe_30_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_18),
		.in_col (out_col_29_19),
		.out_row (out_row_30_19),
		.out_col (out_col_30_19),
		.out_data (out_data_30_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_20;
	wire signed [DATA_WIDTH-1:0] out_col_30_20;
	wire signed [DATA_WIDTH-1:0] out_data_30_20;
	integer_mac_pe mac_pe_30_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_19),
		.in_col (out_col_29_20),
		.out_row (out_row_30_20),
		.out_col (out_col_30_20),
		.out_data (out_data_30_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_21;
	wire signed [DATA_WIDTH-1:0] out_col_30_21;
	wire signed [DATA_WIDTH-1:0] out_data_30_21;
	integer_mac_pe mac_pe_30_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_20),
		.in_col (out_col_29_21),
		.out_row (out_row_30_21),
		.out_col (out_col_30_21),
		.out_data (out_data_30_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_22;
	wire signed [DATA_WIDTH-1:0] out_col_30_22;
	wire signed [DATA_WIDTH-1:0] out_data_30_22;
	integer_mac_pe mac_pe_30_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_21),
		.in_col (out_col_29_22),
		.out_row (out_row_30_22),
		.out_col (out_col_30_22),
		.out_data (out_data_30_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_23;
	wire signed [DATA_WIDTH-1:0] out_col_30_23;
	wire signed [DATA_WIDTH-1:0] out_data_30_23;
	integer_mac_pe mac_pe_30_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_22),
		.in_col (out_col_29_23),
		.out_row (out_row_30_23),
		.out_col (out_col_30_23),
		.out_data (out_data_30_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_24;
	wire signed [DATA_WIDTH-1:0] out_col_30_24;
	wire signed [DATA_WIDTH-1:0] out_data_30_24;
	integer_mac_pe mac_pe_30_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_23),
		.in_col (out_col_29_24),
		.out_row (out_row_30_24),
		.out_col (out_col_30_24),
		.out_data (out_data_30_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_25;
	wire signed [DATA_WIDTH-1:0] out_col_30_25;
	wire signed [DATA_WIDTH-1:0] out_data_30_25;
	integer_mac_pe mac_pe_30_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_24),
		.in_col (out_col_29_25),
		.out_row (out_row_30_25),
		.out_col (out_col_30_25),
		.out_data (out_data_30_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_26;
	wire signed [DATA_WIDTH-1:0] out_col_30_26;
	wire signed [DATA_WIDTH-1:0] out_data_30_26;
	integer_mac_pe mac_pe_30_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_25),
		.in_col (out_col_29_26),
		.out_row (out_row_30_26),
		.out_col (out_col_30_26),
		.out_data (out_data_30_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_27;
	wire signed [DATA_WIDTH-1:0] out_col_30_27;
	wire signed [DATA_WIDTH-1:0] out_data_30_27;
	integer_mac_pe mac_pe_30_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_26),
		.in_col (out_col_29_27),
		.out_row (out_row_30_27),
		.out_col (out_col_30_27),
		.out_data (out_data_30_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_28;
	wire signed [DATA_WIDTH-1:0] out_col_30_28;
	wire signed [DATA_WIDTH-1:0] out_data_30_28;
	integer_mac_pe mac_pe_30_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_27),
		.in_col (out_col_29_28),
		.out_row (out_row_30_28),
		.out_col (out_col_30_28),
		.out_data (out_data_30_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_29;
	wire signed [DATA_WIDTH-1:0] out_col_30_29;
	wire signed [DATA_WIDTH-1:0] out_data_30_29;
	integer_mac_pe mac_pe_30_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_28),
		.in_col (out_col_29_29),
		.out_row (out_row_30_29),
		.out_col (out_col_30_29),
		.out_data (out_data_30_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_30;
	wire signed [DATA_WIDTH-1:0] out_col_30_30;
	wire signed [DATA_WIDTH-1:0] out_data_30_30;
	integer_mac_pe mac_pe_30_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_29),
		.in_col (out_col_29_30),
		.out_row (out_row_30_30),
		.out_col (out_col_30_30),
		.out_data (out_data_30_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_30_31;
	wire signed [DATA_WIDTH-1:0] out_col_30_31;
	wire signed [DATA_WIDTH-1:0] out_data_30_31;
	integer_mac_pe mac_pe_30_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_30_30),
		.in_col (out_col_29_31),
		.out_row (out_row_30_31),
		.out_col (out_col_30_31),
		.out_data (out_data_30_31)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_0;
	wire signed [DATA_WIDTH-1:0] out_col_31_0;
	wire signed [DATA_WIDTH-1:0] out_data_31_0;
	integer_mac_pe mac_pe_31_0 (
		.clk (clk),
		.rstn (rstn),
		.in_row (row_fifo_31_out),
		.in_col (out_col_30_0),
		.out_row (out_row_31_0),
		.out_col (out_col_31_0),
		.out_data (out_data_31_0)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_1;
	wire signed [DATA_WIDTH-1:0] out_col_31_1;
	wire signed [DATA_WIDTH-1:0] out_data_31_1;
	integer_mac_pe mac_pe_31_1 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_0),
		.in_col (out_col_30_1),
		.out_row (out_row_31_1),
		.out_col (out_col_31_1),
		.out_data (out_data_31_1)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_2;
	wire signed [DATA_WIDTH-1:0] out_col_31_2;
	wire signed [DATA_WIDTH-1:0] out_data_31_2;
	integer_mac_pe mac_pe_31_2 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_1),
		.in_col (out_col_30_2),
		.out_row (out_row_31_2),
		.out_col (out_col_31_2),
		.out_data (out_data_31_2)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_3;
	wire signed [DATA_WIDTH-1:0] out_col_31_3;
	wire signed [DATA_WIDTH-1:0] out_data_31_3;
	integer_mac_pe mac_pe_31_3 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_2),
		.in_col (out_col_30_3),
		.out_row (out_row_31_3),
		.out_col (out_col_31_3),
		.out_data (out_data_31_3)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_4;
	wire signed [DATA_WIDTH-1:0] out_col_31_4;
	wire signed [DATA_WIDTH-1:0] out_data_31_4;
	integer_mac_pe mac_pe_31_4 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_3),
		.in_col (out_col_30_4),
		.out_row (out_row_31_4),
		.out_col (out_col_31_4),
		.out_data (out_data_31_4)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_5;
	wire signed [DATA_WIDTH-1:0] out_col_31_5;
	wire signed [DATA_WIDTH-1:0] out_data_31_5;
	integer_mac_pe mac_pe_31_5 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_4),
		.in_col (out_col_30_5),
		.out_row (out_row_31_5),
		.out_col (out_col_31_5),
		.out_data (out_data_31_5)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_6;
	wire signed [DATA_WIDTH-1:0] out_col_31_6;
	wire signed [DATA_WIDTH-1:0] out_data_31_6;
	integer_mac_pe mac_pe_31_6 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_5),
		.in_col (out_col_30_6),
		.out_row (out_row_31_6),
		.out_col (out_col_31_6),
		.out_data (out_data_31_6)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_7;
	wire signed [DATA_WIDTH-1:0] out_col_31_7;
	wire signed [DATA_WIDTH-1:0] out_data_31_7;
	integer_mac_pe mac_pe_31_7 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_6),
		.in_col (out_col_30_7),
		.out_row (out_row_31_7),
		.out_col (out_col_31_7),
		.out_data (out_data_31_7)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_8;
	wire signed [DATA_WIDTH-1:0] out_col_31_8;
	wire signed [DATA_WIDTH-1:0] out_data_31_8;
	integer_mac_pe mac_pe_31_8 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_7),
		.in_col (out_col_30_8),
		.out_row (out_row_31_8),
		.out_col (out_col_31_8),
		.out_data (out_data_31_8)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_9;
	wire signed [DATA_WIDTH-1:0] out_col_31_9;
	wire signed [DATA_WIDTH-1:0] out_data_31_9;
	integer_mac_pe mac_pe_31_9 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_8),
		.in_col (out_col_30_9),
		.out_row (out_row_31_9),
		.out_col (out_col_31_9),
		.out_data (out_data_31_9)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_10;
	wire signed [DATA_WIDTH-1:0] out_col_31_10;
	wire signed [DATA_WIDTH-1:0] out_data_31_10;
	integer_mac_pe mac_pe_31_10 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_9),
		.in_col (out_col_30_10),
		.out_row (out_row_31_10),
		.out_col (out_col_31_10),
		.out_data (out_data_31_10)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_11;
	wire signed [DATA_WIDTH-1:0] out_col_31_11;
	wire signed [DATA_WIDTH-1:0] out_data_31_11;
	integer_mac_pe mac_pe_31_11 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_10),
		.in_col (out_col_30_11),
		.out_row (out_row_31_11),
		.out_col (out_col_31_11),
		.out_data (out_data_31_11)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_12;
	wire signed [DATA_WIDTH-1:0] out_col_31_12;
	wire signed [DATA_WIDTH-1:0] out_data_31_12;
	integer_mac_pe mac_pe_31_12 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_11),
		.in_col (out_col_30_12),
		.out_row (out_row_31_12),
		.out_col (out_col_31_12),
		.out_data (out_data_31_12)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_13;
	wire signed [DATA_WIDTH-1:0] out_col_31_13;
	wire signed [DATA_WIDTH-1:0] out_data_31_13;
	integer_mac_pe mac_pe_31_13 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_12),
		.in_col (out_col_30_13),
		.out_row (out_row_31_13),
		.out_col (out_col_31_13),
		.out_data (out_data_31_13)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_14;
	wire signed [DATA_WIDTH-1:0] out_col_31_14;
	wire signed [DATA_WIDTH-1:0] out_data_31_14;
	integer_mac_pe mac_pe_31_14 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_13),
		.in_col (out_col_30_14),
		.out_row (out_row_31_14),
		.out_col (out_col_31_14),
		.out_data (out_data_31_14)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_15;
	wire signed [DATA_WIDTH-1:0] out_col_31_15;
	wire signed [DATA_WIDTH-1:0] out_data_31_15;
	integer_mac_pe mac_pe_31_15 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_14),
		.in_col (out_col_30_15),
		.out_row (out_row_31_15),
		.out_col (out_col_31_15),
		.out_data (out_data_31_15)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_16;
	wire signed [DATA_WIDTH-1:0] out_col_31_16;
	wire signed [DATA_WIDTH-1:0] out_data_31_16;
	integer_mac_pe mac_pe_31_16 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_15),
		.in_col (out_col_30_16),
		.out_row (out_row_31_16),
		.out_col (out_col_31_16),
		.out_data (out_data_31_16)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_17;
	wire signed [DATA_WIDTH-1:0] out_col_31_17;
	wire signed [DATA_WIDTH-1:0] out_data_31_17;
	integer_mac_pe mac_pe_31_17 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_16),
		.in_col (out_col_30_17),
		.out_row (out_row_31_17),
		.out_col (out_col_31_17),
		.out_data (out_data_31_17)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_18;
	wire signed [DATA_WIDTH-1:0] out_col_31_18;
	wire signed [DATA_WIDTH-1:0] out_data_31_18;
	integer_mac_pe mac_pe_31_18 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_17),
		.in_col (out_col_30_18),
		.out_row (out_row_31_18),
		.out_col (out_col_31_18),
		.out_data (out_data_31_18)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_19;
	wire signed [DATA_WIDTH-1:0] out_col_31_19;
	wire signed [DATA_WIDTH-1:0] out_data_31_19;
	integer_mac_pe mac_pe_31_19 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_18),
		.in_col (out_col_30_19),
		.out_row (out_row_31_19),
		.out_col (out_col_31_19),
		.out_data (out_data_31_19)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_20;
	wire signed [DATA_WIDTH-1:0] out_col_31_20;
	wire signed [DATA_WIDTH-1:0] out_data_31_20;
	integer_mac_pe mac_pe_31_20 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_19),
		.in_col (out_col_30_20),
		.out_row (out_row_31_20),
		.out_col (out_col_31_20),
		.out_data (out_data_31_20)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_21;
	wire signed [DATA_WIDTH-1:0] out_col_31_21;
	wire signed [DATA_WIDTH-1:0] out_data_31_21;
	integer_mac_pe mac_pe_31_21 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_20),
		.in_col (out_col_30_21),
		.out_row (out_row_31_21),
		.out_col (out_col_31_21),
		.out_data (out_data_31_21)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_22;
	wire signed [DATA_WIDTH-1:0] out_col_31_22;
	wire signed [DATA_WIDTH-1:0] out_data_31_22;
	integer_mac_pe mac_pe_31_22 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_21),
		.in_col (out_col_30_22),
		.out_row (out_row_31_22),
		.out_col (out_col_31_22),
		.out_data (out_data_31_22)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_23;
	wire signed [DATA_WIDTH-1:0] out_col_31_23;
	wire signed [DATA_WIDTH-1:0] out_data_31_23;
	integer_mac_pe mac_pe_31_23 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_22),
		.in_col (out_col_30_23),
		.out_row (out_row_31_23),
		.out_col (out_col_31_23),
		.out_data (out_data_31_23)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_24;
	wire signed [DATA_WIDTH-1:0] out_col_31_24;
	wire signed [DATA_WIDTH-1:0] out_data_31_24;
	integer_mac_pe mac_pe_31_24 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_23),
		.in_col (out_col_30_24),
		.out_row (out_row_31_24),
		.out_col (out_col_31_24),
		.out_data (out_data_31_24)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_25;
	wire signed [DATA_WIDTH-1:0] out_col_31_25;
	wire signed [DATA_WIDTH-1:0] out_data_31_25;
	integer_mac_pe mac_pe_31_25 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_24),
		.in_col (out_col_30_25),
		.out_row (out_row_31_25),
		.out_col (out_col_31_25),
		.out_data (out_data_31_25)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_26;
	wire signed [DATA_WIDTH-1:0] out_col_31_26;
	wire signed [DATA_WIDTH-1:0] out_data_31_26;
	integer_mac_pe mac_pe_31_26 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_25),
		.in_col (out_col_30_26),
		.out_row (out_row_31_26),
		.out_col (out_col_31_26),
		.out_data (out_data_31_26)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_27;
	wire signed [DATA_WIDTH-1:0] out_col_31_27;
	wire signed [DATA_WIDTH-1:0] out_data_31_27;
	integer_mac_pe mac_pe_31_27 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_26),
		.in_col (out_col_30_27),
		.out_row (out_row_31_27),
		.out_col (out_col_31_27),
		.out_data (out_data_31_27)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_28;
	wire signed [DATA_WIDTH-1:0] out_col_31_28;
	wire signed [DATA_WIDTH-1:0] out_data_31_28;
	integer_mac_pe mac_pe_31_28 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_27),
		.in_col (out_col_30_28),
		.out_row (out_row_31_28),
		.out_col (out_col_31_28),
		.out_data (out_data_31_28)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_29;
	wire signed [DATA_WIDTH-1:0] out_col_31_29;
	wire signed [DATA_WIDTH-1:0] out_data_31_29;
	integer_mac_pe mac_pe_31_29 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_28),
		.in_col (out_col_30_29),
		.out_row (out_row_31_29),
		.out_col (out_col_31_29),
		.out_data (out_data_31_29)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_30;
	wire signed [DATA_WIDTH-1:0] out_col_31_30;
	wire signed [DATA_WIDTH-1:0] out_data_31_30;
	integer_mac_pe mac_pe_31_30 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_29),
		.in_col (out_col_30_30),
		.out_row (out_row_31_30),
		.out_col (out_col_31_30),
		.out_data (out_data_31_30)
	);
	wire signed [DATA_WIDTH-1:0] out_row_31_31;
	wire signed [DATA_WIDTH-1:0] out_col_31_31;
	wire signed [DATA_WIDTH-1:0] out_data_31_31;
	integer_mac_pe mac_pe_31_31 (
		.clk (clk),
		.rstn (rstn),
		.in_row (out_row_31_30),
		.in_col (out_col_30_31),
		.out_row (out_row_31_31),
		.out_col (out_col_31_31),
		.out_data (out_data_31_31)
	);
	mux_1024_to_1  mux (
		.select (out_select),
		.in_data_0_0 (out_data_0_0),
		.in_data_0_1 (out_data_0_1),
		.in_data_0_2 (out_data_0_2),
		.in_data_0_3 (out_data_0_3),
		.in_data_0_4 (out_data_0_4),
		.in_data_0_5 (out_data_0_5),
		.in_data_0_6 (out_data_0_6),
		.in_data_0_7 (out_data_0_7),
		.in_data_0_8 (out_data_0_8),
		.in_data_0_9 (out_data_0_9),
		.in_data_0_10 (out_data_0_10),
		.in_data_0_11 (out_data_0_11),
		.in_data_0_12 (out_data_0_12),
		.in_data_0_13 (out_data_0_13),
		.in_data_0_14 (out_data_0_14),
		.in_data_0_15 (out_data_0_15),
		.in_data_0_16 (out_data_0_16),
		.in_data_0_17 (out_data_0_17),
		.in_data_0_18 (out_data_0_18),
		.in_data_0_19 (out_data_0_19),
		.in_data_0_20 (out_data_0_20),
		.in_data_0_21 (out_data_0_21),
		.in_data_0_22 (out_data_0_22),
		.in_data_0_23 (out_data_0_23),
		.in_data_0_24 (out_data_0_24),
		.in_data_0_25 (out_data_0_25),
		.in_data_0_26 (out_data_0_26),
		.in_data_0_27 (out_data_0_27),
		.in_data_0_28 (out_data_0_28),
		.in_data_0_29 (out_data_0_29),
		.in_data_0_30 (out_data_0_30),
		.in_data_0_31 (out_data_0_31),
		.in_data_1_0 (out_data_1_0),
		.in_data_1_1 (out_data_1_1),
		.in_data_1_2 (out_data_1_2),
		.in_data_1_3 (out_data_1_3),
		.in_data_1_4 (out_data_1_4),
		.in_data_1_5 (out_data_1_5),
		.in_data_1_6 (out_data_1_6),
		.in_data_1_7 (out_data_1_7),
		.in_data_1_8 (out_data_1_8),
		.in_data_1_9 (out_data_1_9),
		.in_data_1_10 (out_data_1_10),
		.in_data_1_11 (out_data_1_11),
		.in_data_1_12 (out_data_1_12),
		.in_data_1_13 (out_data_1_13),
		.in_data_1_14 (out_data_1_14),
		.in_data_1_15 (out_data_1_15),
		.in_data_1_16 (out_data_1_16),
		.in_data_1_17 (out_data_1_17),
		.in_data_1_18 (out_data_1_18),
		.in_data_1_19 (out_data_1_19),
		.in_data_1_20 (out_data_1_20),
		.in_data_1_21 (out_data_1_21),
		.in_data_1_22 (out_data_1_22),
		.in_data_1_23 (out_data_1_23),
		.in_data_1_24 (out_data_1_24),
		.in_data_1_25 (out_data_1_25),
		.in_data_1_26 (out_data_1_26),
		.in_data_1_27 (out_data_1_27),
		.in_data_1_28 (out_data_1_28),
		.in_data_1_29 (out_data_1_29),
		.in_data_1_30 (out_data_1_30),
		.in_data_1_31 (out_data_1_31),
		.in_data_2_0 (out_data_2_0),
		.in_data_2_1 (out_data_2_1),
		.in_data_2_2 (out_data_2_2),
		.in_data_2_3 (out_data_2_3),
		.in_data_2_4 (out_data_2_4),
		.in_data_2_5 (out_data_2_5),
		.in_data_2_6 (out_data_2_6),
		.in_data_2_7 (out_data_2_7),
		.in_data_2_8 (out_data_2_8),
		.in_data_2_9 (out_data_2_9),
		.in_data_2_10 (out_data_2_10),
		.in_data_2_11 (out_data_2_11),
		.in_data_2_12 (out_data_2_12),
		.in_data_2_13 (out_data_2_13),
		.in_data_2_14 (out_data_2_14),
		.in_data_2_15 (out_data_2_15),
		.in_data_2_16 (out_data_2_16),
		.in_data_2_17 (out_data_2_17),
		.in_data_2_18 (out_data_2_18),
		.in_data_2_19 (out_data_2_19),
		.in_data_2_20 (out_data_2_20),
		.in_data_2_21 (out_data_2_21),
		.in_data_2_22 (out_data_2_22),
		.in_data_2_23 (out_data_2_23),
		.in_data_2_24 (out_data_2_24),
		.in_data_2_25 (out_data_2_25),
		.in_data_2_26 (out_data_2_26),
		.in_data_2_27 (out_data_2_27),
		.in_data_2_28 (out_data_2_28),
		.in_data_2_29 (out_data_2_29),
		.in_data_2_30 (out_data_2_30),
		.in_data_2_31 (out_data_2_31),
		.in_data_3_0 (out_data_3_0),
		.in_data_3_1 (out_data_3_1),
		.in_data_3_2 (out_data_3_2),
		.in_data_3_3 (out_data_3_3),
		.in_data_3_4 (out_data_3_4),
		.in_data_3_5 (out_data_3_5),
		.in_data_3_6 (out_data_3_6),
		.in_data_3_7 (out_data_3_7),
		.in_data_3_8 (out_data_3_8),
		.in_data_3_9 (out_data_3_9),
		.in_data_3_10 (out_data_3_10),
		.in_data_3_11 (out_data_3_11),
		.in_data_3_12 (out_data_3_12),
		.in_data_3_13 (out_data_3_13),
		.in_data_3_14 (out_data_3_14),
		.in_data_3_15 (out_data_3_15),
		.in_data_3_16 (out_data_3_16),
		.in_data_3_17 (out_data_3_17),
		.in_data_3_18 (out_data_3_18),
		.in_data_3_19 (out_data_3_19),
		.in_data_3_20 (out_data_3_20),
		.in_data_3_21 (out_data_3_21),
		.in_data_3_22 (out_data_3_22),
		.in_data_3_23 (out_data_3_23),
		.in_data_3_24 (out_data_3_24),
		.in_data_3_25 (out_data_3_25),
		.in_data_3_26 (out_data_3_26),
		.in_data_3_27 (out_data_3_27),
		.in_data_3_28 (out_data_3_28),
		.in_data_3_29 (out_data_3_29),
		.in_data_3_30 (out_data_3_30),
		.in_data_3_31 (out_data_3_31),
		.in_data_4_0 (out_data_4_0),
		.in_data_4_1 (out_data_4_1),
		.in_data_4_2 (out_data_4_2),
		.in_data_4_3 (out_data_4_3),
		.in_data_4_4 (out_data_4_4),
		.in_data_4_5 (out_data_4_5),
		.in_data_4_6 (out_data_4_6),
		.in_data_4_7 (out_data_4_7),
		.in_data_4_8 (out_data_4_8),
		.in_data_4_9 (out_data_4_9),
		.in_data_4_10 (out_data_4_10),
		.in_data_4_11 (out_data_4_11),
		.in_data_4_12 (out_data_4_12),
		.in_data_4_13 (out_data_4_13),
		.in_data_4_14 (out_data_4_14),
		.in_data_4_15 (out_data_4_15),
		.in_data_4_16 (out_data_4_16),
		.in_data_4_17 (out_data_4_17),
		.in_data_4_18 (out_data_4_18),
		.in_data_4_19 (out_data_4_19),
		.in_data_4_20 (out_data_4_20),
		.in_data_4_21 (out_data_4_21),
		.in_data_4_22 (out_data_4_22),
		.in_data_4_23 (out_data_4_23),
		.in_data_4_24 (out_data_4_24),
		.in_data_4_25 (out_data_4_25),
		.in_data_4_26 (out_data_4_26),
		.in_data_4_27 (out_data_4_27),
		.in_data_4_28 (out_data_4_28),
		.in_data_4_29 (out_data_4_29),
		.in_data_4_30 (out_data_4_30),
		.in_data_4_31 (out_data_4_31),
		.in_data_5_0 (out_data_5_0),
		.in_data_5_1 (out_data_5_1),
		.in_data_5_2 (out_data_5_2),
		.in_data_5_3 (out_data_5_3),
		.in_data_5_4 (out_data_5_4),
		.in_data_5_5 (out_data_5_5),
		.in_data_5_6 (out_data_5_6),
		.in_data_5_7 (out_data_5_7),
		.in_data_5_8 (out_data_5_8),
		.in_data_5_9 (out_data_5_9),
		.in_data_5_10 (out_data_5_10),
		.in_data_5_11 (out_data_5_11),
		.in_data_5_12 (out_data_5_12),
		.in_data_5_13 (out_data_5_13),
		.in_data_5_14 (out_data_5_14),
		.in_data_5_15 (out_data_5_15),
		.in_data_5_16 (out_data_5_16),
		.in_data_5_17 (out_data_5_17),
		.in_data_5_18 (out_data_5_18),
		.in_data_5_19 (out_data_5_19),
		.in_data_5_20 (out_data_5_20),
		.in_data_5_21 (out_data_5_21),
		.in_data_5_22 (out_data_5_22),
		.in_data_5_23 (out_data_5_23),
		.in_data_5_24 (out_data_5_24),
		.in_data_5_25 (out_data_5_25),
		.in_data_5_26 (out_data_5_26),
		.in_data_5_27 (out_data_5_27),
		.in_data_5_28 (out_data_5_28),
		.in_data_5_29 (out_data_5_29),
		.in_data_5_30 (out_data_5_30),
		.in_data_5_31 (out_data_5_31),
		.in_data_6_0 (out_data_6_0),
		.in_data_6_1 (out_data_6_1),
		.in_data_6_2 (out_data_6_2),
		.in_data_6_3 (out_data_6_3),
		.in_data_6_4 (out_data_6_4),
		.in_data_6_5 (out_data_6_5),
		.in_data_6_6 (out_data_6_6),
		.in_data_6_7 (out_data_6_7),
		.in_data_6_8 (out_data_6_8),
		.in_data_6_9 (out_data_6_9),
		.in_data_6_10 (out_data_6_10),
		.in_data_6_11 (out_data_6_11),
		.in_data_6_12 (out_data_6_12),
		.in_data_6_13 (out_data_6_13),
		.in_data_6_14 (out_data_6_14),
		.in_data_6_15 (out_data_6_15),
		.in_data_6_16 (out_data_6_16),
		.in_data_6_17 (out_data_6_17),
		.in_data_6_18 (out_data_6_18),
		.in_data_6_19 (out_data_6_19),
		.in_data_6_20 (out_data_6_20),
		.in_data_6_21 (out_data_6_21),
		.in_data_6_22 (out_data_6_22),
		.in_data_6_23 (out_data_6_23),
		.in_data_6_24 (out_data_6_24),
		.in_data_6_25 (out_data_6_25),
		.in_data_6_26 (out_data_6_26),
		.in_data_6_27 (out_data_6_27),
		.in_data_6_28 (out_data_6_28),
		.in_data_6_29 (out_data_6_29),
		.in_data_6_30 (out_data_6_30),
		.in_data_6_31 (out_data_6_31),
		.in_data_7_0 (out_data_7_0),
		.in_data_7_1 (out_data_7_1),
		.in_data_7_2 (out_data_7_2),
		.in_data_7_3 (out_data_7_3),
		.in_data_7_4 (out_data_7_4),
		.in_data_7_5 (out_data_7_5),
		.in_data_7_6 (out_data_7_6),
		.in_data_7_7 (out_data_7_7),
		.in_data_7_8 (out_data_7_8),
		.in_data_7_9 (out_data_7_9),
		.in_data_7_10 (out_data_7_10),
		.in_data_7_11 (out_data_7_11),
		.in_data_7_12 (out_data_7_12),
		.in_data_7_13 (out_data_7_13),
		.in_data_7_14 (out_data_7_14),
		.in_data_7_15 (out_data_7_15),
		.in_data_7_16 (out_data_7_16),
		.in_data_7_17 (out_data_7_17),
		.in_data_7_18 (out_data_7_18),
		.in_data_7_19 (out_data_7_19),
		.in_data_7_20 (out_data_7_20),
		.in_data_7_21 (out_data_7_21),
		.in_data_7_22 (out_data_7_22),
		.in_data_7_23 (out_data_7_23),
		.in_data_7_24 (out_data_7_24),
		.in_data_7_25 (out_data_7_25),
		.in_data_7_26 (out_data_7_26),
		.in_data_7_27 (out_data_7_27),
		.in_data_7_28 (out_data_7_28),
		.in_data_7_29 (out_data_7_29),
		.in_data_7_30 (out_data_7_30),
		.in_data_7_31 (out_data_7_31),
		.in_data_8_0 (out_data_8_0),
		.in_data_8_1 (out_data_8_1),
		.in_data_8_2 (out_data_8_2),
		.in_data_8_3 (out_data_8_3),
		.in_data_8_4 (out_data_8_4),
		.in_data_8_5 (out_data_8_5),
		.in_data_8_6 (out_data_8_6),
		.in_data_8_7 (out_data_8_7),
		.in_data_8_8 (out_data_8_8),
		.in_data_8_9 (out_data_8_9),
		.in_data_8_10 (out_data_8_10),
		.in_data_8_11 (out_data_8_11),
		.in_data_8_12 (out_data_8_12),
		.in_data_8_13 (out_data_8_13),
		.in_data_8_14 (out_data_8_14),
		.in_data_8_15 (out_data_8_15),
		.in_data_8_16 (out_data_8_16),
		.in_data_8_17 (out_data_8_17),
		.in_data_8_18 (out_data_8_18),
		.in_data_8_19 (out_data_8_19),
		.in_data_8_20 (out_data_8_20),
		.in_data_8_21 (out_data_8_21),
		.in_data_8_22 (out_data_8_22),
		.in_data_8_23 (out_data_8_23),
		.in_data_8_24 (out_data_8_24),
		.in_data_8_25 (out_data_8_25),
		.in_data_8_26 (out_data_8_26),
		.in_data_8_27 (out_data_8_27),
		.in_data_8_28 (out_data_8_28),
		.in_data_8_29 (out_data_8_29),
		.in_data_8_30 (out_data_8_30),
		.in_data_8_31 (out_data_8_31),
		.in_data_9_0 (out_data_9_0),
		.in_data_9_1 (out_data_9_1),
		.in_data_9_2 (out_data_9_2),
		.in_data_9_3 (out_data_9_3),
		.in_data_9_4 (out_data_9_4),
		.in_data_9_5 (out_data_9_5),
		.in_data_9_6 (out_data_9_6),
		.in_data_9_7 (out_data_9_7),
		.in_data_9_8 (out_data_9_8),
		.in_data_9_9 (out_data_9_9),
		.in_data_9_10 (out_data_9_10),
		.in_data_9_11 (out_data_9_11),
		.in_data_9_12 (out_data_9_12),
		.in_data_9_13 (out_data_9_13),
		.in_data_9_14 (out_data_9_14),
		.in_data_9_15 (out_data_9_15),
		.in_data_9_16 (out_data_9_16),
		.in_data_9_17 (out_data_9_17),
		.in_data_9_18 (out_data_9_18),
		.in_data_9_19 (out_data_9_19),
		.in_data_9_20 (out_data_9_20),
		.in_data_9_21 (out_data_9_21),
		.in_data_9_22 (out_data_9_22),
		.in_data_9_23 (out_data_9_23),
		.in_data_9_24 (out_data_9_24),
		.in_data_9_25 (out_data_9_25),
		.in_data_9_26 (out_data_9_26),
		.in_data_9_27 (out_data_9_27),
		.in_data_9_28 (out_data_9_28),
		.in_data_9_29 (out_data_9_29),
		.in_data_9_30 (out_data_9_30),
		.in_data_9_31 (out_data_9_31),
		.in_data_10_0 (out_data_10_0),
		.in_data_10_1 (out_data_10_1),
		.in_data_10_2 (out_data_10_2),
		.in_data_10_3 (out_data_10_3),
		.in_data_10_4 (out_data_10_4),
		.in_data_10_5 (out_data_10_5),
		.in_data_10_6 (out_data_10_6),
		.in_data_10_7 (out_data_10_7),
		.in_data_10_8 (out_data_10_8),
		.in_data_10_9 (out_data_10_9),
		.in_data_10_10 (out_data_10_10),
		.in_data_10_11 (out_data_10_11),
		.in_data_10_12 (out_data_10_12),
		.in_data_10_13 (out_data_10_13),
		.in_data_10_14 (out_data_10_14),
		.in_data_10_15 (out_data_10_15),
		.in_data_10_16 (out_data_10_16),
		.in_data_10_17 (out_data_10_17),
		.in_data_10_18 (out_data_10_18),
		.in_data_10_19 (out_data_10_19),
		.in_data_10_20 (out_data_10_20),
		.in_data_10_21 (out_data_10_21),
		.in_data_10_22 (out_data_10_22),
		.in_data_10_23 (out_data_10_23),
		.in_data_10_24 (out_data_10_24),
		.in_data_10_25 (out_data_10_25),
		.in_data_10_26 (out_data_10_26),
		.in_data_10_27 (out_data_10_27),
		.in_data_10_28 (out_data_10_28),
		.in_data_10_29 (out_data_10_29),
		.in_data_10_30 (out_data_10_30),
		.in_data_10_31 (out_data_10_31),
		.in_data_11_0 (out_data_11_0),
		.in_data_11_1 (out_data_11_1),
		.in_data_11_2 (out_data_11_2),
		.in_data_11_3 (out_data_11_3),
		.in_data_11_4 (out_data_11_4),
		.in_data_11_5 (out_data_11_5),
		.in_data_11_6 (out_data_11_6),
		.in_data_11_7 (out_data_11_7),
		.in_data_11_8 (out_data_11_8),
		.in_data_11_9 (out_data_11_9),
		.in_data_11_10 (out_data_11_10),
		.in_data_11_11 (out_data_11_11),
		.in_data_11_12 (out_data_11_12),
		.in_data_11_13 (out_data_11_13),
		.in_data_11_14 (out_data_11_14),
		.in_data_11_15 (out_data_11_15),
		.in_data_11_16 (out_data_11_16),
		.in_data_11_17 (out_data_11_17),
		.in_data_11_18 (out_data_11_18),
		.in_data_11_19 (out_data_11_19),
		.in_data_11_20 (out_data_11_20),
		.in_data_11_21 (out_data_11_21),
		.in_data_11_22 (out_data_11_22),
		.in_data_11_23 (out_data_11_23),
		.in_data_11_24 (out_data_11_24),
		.in_data_11_25 (out_data_11_25),
		.in_data_11_26 (out_data_11_26),
		.in_data_11_27 (out_data_11_27),
		.in_data_11_28 (out_data_11_28),
		.in_data_11_29 (out_data_11_29),
		.in_data_11_30 (out_data_11_30),
		.in_data_11_31 (out_data_11_31),
		.in_data_12_0 (out_data_12_0),
		.in_data_12_1 (out_data_12_1),
		.in_data_12_2 (out_data_12_2),
		.in_data_12_3 (out_data_12_3),
		.in_data_12_4 (out_data_12_4),
		.in_data_12_5 (out_data_12_5),
		.in_data_12_6 (out_data_12_6),
		.in_data_12_7 (out_data_12_7),
		.in_data_12_8 (out_data_12_8),
		.in_data_12_9 (out_data_12_9),
		.in_data_12_10 (out_data_12_10),
		.in_data_12_11 (out_data_12_11),
		.in_data_12_12 (out_data_12_12),
		.in_data_12_13 (out_data_12_13),
		.in_data_12_14 (out_data_12_14),
		.in_data_12_15 (out_data_12_15),
		.in_data_12_16 (out_data_12_16),
		.in_data_12_17 (out_data_12_17),
		.in_data_12_18 (out_data_12_18),
		.in_data_12_19 (out_data_12_19),
		.in_data_12_20 (out_data_12_20),
		.in_data_12_21 (out_data_12_21),
		.in_data_12_22 (out_data_12_22),
		.in_data_12_23 (out_data_12_23),
		.in_data_12_24 (out_data_12_24),
		.in_data_12_25 (out_data_12_25),
		.in_data_12_26 (out_data_12_26),
		.in_data_12_27 (out_data_12_27),
		.in_data_12_28 (out_data_12_28),
		.in_data_12_29 (out_data_12_29),
		.in_data_12_30 (out_data_12_30),
		.in_data_12_31 (out_data_12_31),
		.in_data_13_0 (out_data_13_0),
		.in_data_13_1 (out_data_13_1),
		.in_data_13_2 (out_data_13_2),
		.in_data_13_3 (out_data_13_3),
		.in_data_13_4 (out_data_13_4),
		.in_data_13_5 (out_data_13_5),
		.in_data_13_6 (out_data_13_6),
		.in_data_13_7 (out_data_13_7),
		.in_data_13_8 (out_data_13_8),
		.in_data_13_9 (out_data_13_9),
		.in_data_13_10 (out_data_13_10),
		.in_data_13_11 (out_data_13_11),
		.in_data_13_12 (out_data_13_12),
		.in_data_13_13 (out_data_13_13),
		.in_data_13_14 (out_data_13_14),
		.in_data_13_15 (out_data_13_15),
		.in_data_13_16 (out_data_13_16),
		.in_data_13_17 (out_data_13_17),
		.in_data_13_18 (out_data_13_18),
		.in_data_13_19 (out_data_13_19),
		.in_data_13_20 (out_data_13_20),
		.in_data_13_21 (out_data_13_21),
		.in_data_13_22 (out_data_13_22),
		.in_data_13_23 (out_data_13_23),
		.in_data_13_24 (out_data_13_24),
		.in_data_13_25 (out_data_13_25),
		.in_data_13_26 (out_data_13_26),
		.in_data_13_27 (out_data_13_27),
		.in_data_13_28 (out_data_13_28),
		.in_data_13_29 (out_data_13_29),
		.in_data_13_30 (out_data_13_30),
		.in_data_13_31 (out_data_13_31),
		.in_data_14_0 (out_data_14_0),
		.in_data_14_1 (out_data_14_1),
		.in_data_14_2 (out_data_14_2),
		.in_data_14_3 (out_data_14_3),
		.in_data_14_4 (out_data_14_4),
		.in_data_14_5 (out_data_14_5),
		.in_data_14_6 (out_data_14_6),
		.in_data_14_7 (out_data_14_7),
		.in_data_14_8 (out_data_14_8),
		.in_data_14_9 (out_data_14_9),
		.in_data_14_10 (out_data_14_10),
		.in_data_14_11 (out_data_14_11),
		.in_data_14_12 (out_data_14_12),
		.in_data_14_13 (out_data_14_13),
		.in_data_14_14 (out_data_14_14),
		.in_data_14_15 (out_data_14_15),
		.in_data_14_16 (out_data_14_16),
		.in_data_14_17 (out_data_14_17),
		.in_data_14_18 (out_data_14_18),
		.in_data_14_19 (out_data_14_19),
		.in_data_14_20 (out_data_14_20),
		.in_data_14_21 (out_data_14_21),
		.in_data_14_22 (out_data_14_22),
		.in_data_14_23 (out_data_14_23),
		.in_data_14_24 (out_data_14_24),
		.in_data_14_25 (out_data_14_25),
		.in_data_14_26 (out_data_14_26),
		.in_data_14_27 (out_data_14_27),
		.in_data_14_28 (out_data_14_28),
		.in_data_14_29 (out_data_14_29),
		.in_data_14_30 (out_data_14_30),
		.in_data_14_31 (out_data_14_31),
		.in_data_15_0 (out_data_15_0),
		.in_data_15_1 (out_data_15_1),
		.in_data_15_2 (out_data_15_2),
		.in_data_15_3 (out_data_15_3),
		.in_data_15_4 (out_data_15_4),
		.in_data_15_5 (out_data_15_5),
		.in_data_15_6 (out_data_15_6),
		.in_data_15_7 (out_data_15_7),
		.in_data_15_8 (out_data_15_8),
		.in_data_15_9 (out_data_15_9),
		.in_data_15_10 (out_data_15_10),
		.in_data_15_11 (out_data_15_11),
		.in_data_15_12 (out_data_15_12),
		.in_data_15_13 (out_data_15_13),
		.in_data_15_14 (out_data_15_14),
		.in_data_15_15 (out_data_15_15),
		.in_data_15_16 (out_data_15_16),
		.in_data_15_17 (out_data_15_17),
		.in_data_15_18 (out_data_15_18),
		.in_data_15_19 (out_data_15_19),
		.in_data_15_20 (out_data_15_20),
		.in_data_15_21 (out_data_15_21),
		.in_data_15_22 (out_data_15_22),
		.in_data_15_23 (out_data_15_23),
		.in_data_15_24 (out_data_15_24),
		.in_data_15_25 (out_data_15_25),
		.in_data_15_26 (out_data_15_26),
		.in_data_15_27 (out_data_15_27),
		.in_data_15_28 (out_data_15_28),
		.in_data_15_29 (out_data_15_29),
		.in_data_15_30 (out_data_15_30),
		.in_data_15_31 (out_data_15_31),
		.in_data_16_0 (out_data_16_0),
		.in_data_16_1 (out_data_16_1),
		.in_data_16_2 (out_data_16_2),
		.in_data_16_3 (out_data_16_3),
		.in_data_16_4 (out_data_16_4),
		.in_data_16_5 (out_data_16_5),
		.in_data_16_6 (out_data_16_6),
		.in_data_16_7 (out_data_16_7),
		.in_data_16_8 (out_data_16_8),
		.in_data_16_9 (out_data_16_9),
		.in_data_16_10 (out_data_16_10),
		.in_data_16_11 (out_data_16_11),
		.in_data_16_12 (out_data_16_12),
		.in_data_16_13 (out_data_16_13),
		.in_data_16_14 (out_data_16_14),
		.in_data_16_15 (out_data_16_15),
		.in_data_16_16 (out_data_16_16),
		.in_data_16_17 (out_data_16_17),
		.in_data_16_18 (out_data_16_18),
		.in_data_16_19 (out_data_16_19),
		.in_data_16_20 (out_data_16_20),
		.in_data_16_21 (out_data_16_21),
		.in_data_16_22 (out_data_16_22),
		.in_data_16_23 (out_data_16_23),
		.in_data_16_24 (out_data_16_24),
		.in_data_16_25 (out_data_16_25),
		.in_data_16_26 (out_data_16_26),
		.in_data_16_27 (out_data_16_27),
		.in_data_16_28 (out_data_16_28),
		.in_data_16_29 (out_data_16_29),
		.in_data_16_30 (out_data_16_30),
		.in_data_16_31 (out_data_16_31),
		.in_data_17_0 (out_data_17_0),
		.in_data_17_1 (out_data_17_1),
		.in_data_17_2 (out_data_17_2),
		.in_data_17_3 (out_data_17_3),
		.in_data_17_4 (out_data_17_4),
		.in_data_17_5 (out_data_17_5),
		.in_data_17_6 (out_data_17_6),
		.in_data_17_7 (out_data_17_7),
		.in_data_17_8 (out_data_17_8),
		.in_data_17_9 (out_data_17_9),
		.in_data_17_10 (out_data_17_10),
		.in_data_17_11 (out_data_17_11),
		.in_data_17_12 (out_data_17_12),
		.in_data_17_13 (out_data_17_13),
		.in_data_17_14 (out_data_17_14),
		.in_data_17_15 (out_data_17_15),
		.in_data_17_16 (out_data_17_16),
		.in_data_17_17 (out_data_17_17),
		.in_data_17_18 (out_data_17_18),
		.in_data_17_19 (out_data_17_19),
		.in_data_17_20 (out_data_17_20),
		.in_data_17_21 (out_data_17_21),
		.in_data_17_22 (out_data_17_22),
		.in_data_17_23 (out_data_17_23),
		.in_data_17_24 (out_data_17_24),
		.in_data_17_25 (out_data_17_25),
		.in_data_17_26 (out_data_17_26),
		.in_data_17_27 (out_data_17_27),
		.in_data_17_28 (out_data_17_28),
		.in_data_17_29 (out_data_17_29),
		.in_data_17_30 (out_data_17_30),
		.in_data_17_31 (out_data_17_31),
		.in_data_18_0 (out_data_18_0),
		.in_data_18_1 (out_data_18_1),
		.in_data_18_2 (out_data_18_2),
		.in_data_18_3 (out_data_18_3),
		.in_data_18_4 (out_data_18_4),
		.in_data_18_5 (out_data_18_5),
		.in_data_18_6 (out_data_18_6),
		.in_data_18_7 (out_data_18_7),
		.in_data_18_8 (out_data_18_8),
		.in_data_18_9 (out_data_18_9),
		.in_data_18_10 (out_data_18_10),
		.in_data_18_11 (out_data_18_11),
		.in_data_18_12 (out_data_18_12),
		.in_data_18_13 (out_data_18_13),
		.in_data_18_14 (out_data_18_14),
		.in_data_18_15 (out_data_18_15),
		.in_data_18_16 (out_data_18_16),
		.in_data_18_17 (out_data_18_17),
		.in_data_18_18 (out_data_18_18),
		.in_data_18_19 (out_data_18_19),
		.in_data_18_20 (out_data_18_20),
		.in_data_18_21 (out_data_18_21),
		.in_data_18_22 (out_data_18_22),
		.in_data_18_23 (out_data_18_23),
		.in_data_18_24 (out_data_18_24),
		.in_data_18_25 (out_data_18_25),
		.in_data_18_26 (out_data_18_26),
		.in_data_18_27 (out_data_18_27),
		.in_data_18_28 (out_data_18_28),
		.in_data_18_29 (out_data_18_29),
		.in_data_18_30 (out_data_18_30),
		.in_data_18_31 (out_data_18_31),
		.in_data_19_0 (out_data_19_0),
		.in_data_19_1 (out_data_19_1),
		.in_data_19_2 (out_data_19_2),
		.in_data_19_3 (out_data_19_3),
		.in_data_19_4 (out_data_19_4),
		.in_data_19_5 (out_data_19_5),
		.in_data_19_6 (out_data_19_6),
		.in_data_19_7 (out_data_19_7),
		.in_data_19_8 (out_data_19_8),
		.in_data_19_9 (out_data_19_9),
		.in_data_19_10 (out_data_19_10),
		.in_data_19_11 (out_data_19_11),
		.in_data_19_12 (out_data_19_12),
		.in_data_19_13 (out_data_19_13),
		.in_data_19_14 (out_data_19_14),
		.in_data_19_15 (out_data_19_15),
		.in_data_19_16 (out_data_19_16),
		.in_data_19_17 (out_data_19_17),
		.in_data_19_18 (out_data_19_18),
		.in_data_19_19 (out_data_19_19),
		.in_data_19_20 (out_data_19_20),
		.in_data_19_21 (out_data_19_21),
		.in_data_19_22 (out_data_19_22),
		.in_data_19_23 (out_data_19_23),
		.in_data_19_24 (out_data_19_24),
		.in_data_19_25 (out_data_19_25),
		.in_data_19_26 (out_data_19_26),
		.in_data_19_27 (out_data_19_27),
		.in_data_19_28 (out_data_19_28),
		.in_data_19_29 (out_data_19_29),
		.in_data_19_30 (out_data_19_30),
		.in_data_19_31 (out_data_19_31),
		.in_data_20_0 (out_data_20_0),
		.in_data_20_1 (out_data_20_1),
		.in_data_20_2 (out_data_20_2),
		.in_data_20_3 (out_data_20_3),
		.in_data_20_4 (out_data_20_4),
		.in_data_20_5 (out_data_20_5),
		.in_data_20_6 (out_data_20_6),
		.in_data_20_7 (out_data_20_7),
		.in_data_20_8 (out_data_20_8),
		.in_data_20_9 (out_data_20_9),
		.in_data_20_10 (out_data_20_10),
		.in_data_20_11 (out_data_20_11),
		.in_data_20_12 (out_data_20_12),
		.in_data_20_13 (out_data_20_13),
		.in_data_20_14 (out_data_20_14),
		.in_data_20_15 (out_data_20_15),
		.in_data_20_16 (out_data_20_16),
		.in_data_20_17 (out_data_20_17),
		.in_data_20_18 (out_data_20_18),
		.in_data_20_19 (out_data_20_19),
		.in_data_20_20 (out_data_20_20),
		.in_data_20_21 (out_data_20_21),
		.in_data_20_22 (out_data_20_22),
		.in_data_20_23 (out_data_20_23),
		.in_data_20_24 (out_data_20_24),
		.in_data_20_25 (out_data_20_25),
		.in_data_20_26 (out_data_20_26),
		.in_data_20_27 (out_data_20_27),
		.in_data_20_28 (out_data_20_28),
		.in_data_20_29 (out_data_20_29),
		.in_data_20_30 (out_data_20_30),
		.in_data_20_31 (out_data_20_31),
		.in_data_21_0 (out_data_21_0),
		.in_data_21_1 (out_data_21_1),
		.in_data_21_2 (out_data_21_2),
		.in_data_21_3 (out_data_21_3),
		.in_data_21_4 (out_data_21_4),
		.in_data_21_5 (out_data_21_5),
		.in_data_21_6 (out_data_21_6),
		.in_data_21_7 (out_data_21_7),
		.in_data_21_8 (out_data_21_8),
		.in_data_21_9 (out_data_21_9),
		.in_data_21_10 (out_data_21_10),
		.in_data_21_11 (out_data_21_11),
		.in_data_21_12 (out_data_21_12),
		.in_data_21_13 (out_data_21_13),
		.in_data_21_14 (out_data_21_14),
		.in_data_21_15 (out_data_21_15),
		.in_data_21_16 (out_data_21_16),
		.in_data_21_17 (out_data_21_17),
		.in_data_21_18 (out_data_21_18),
		.in_data_21_19 (out_data_21_19),
		.in_data_21_20 (out_data_21_20),
		.in_data_21_21 (out_data_21_21),
		.in_data_21_22 (out_data_21_22),
		.in_data_21_23 (out_data_21_23),
		.in_data_21_24 (out_data_21_24),
		.in_data_21_25 (out_data_21_25),
		.in_data_21_26 (out_data_21_26),
		.in_data_21_27 (out_data_21_27),
		.in_data_21_28 (out_data_21_28),
		.in_data_21_29 (out_data_21_29),
		.in_data_21_30 (out_data_21_30),
		.in_data_21_31 (out_data_21_31),
		.in_data_22_0 (out_data_22_0),
		.in_data_22_1 (out_data_22_1),
		.in_data_22_2 (out_data_22_2),
		.in_data_22_3 (out_data_22_3),
		.in_data_22_4 (out_data_22_4),
		.in_data_22_5 (out_data_22_5),
		.in_data_22_6 (out_data_22_6),
		.in_data_22_7 (out_data_22_7),
		.in_data_22_8 (out_data_22_8),
		.in_data_22_9 (out_data_22_9),
		.in_data_22_10 (out_data_22_10),
		.in_data_22_11 (out_data_22_11),
		.in_data_22_12 (out_data_22_12),
		.in_data_22_13 (out_data_22_13),
		.in_data_22_14 (out_data_22_14),
		.in_data_22_15 (out_data_22_15),
		.in_data_22_16 (out_data_22_16),
		.in_data_22_17 (out_data_22_17),
		.in_data_22_18 (out_data_22_18),
		.in_data_22_19 (out_data_22_19),
		.in_data_22_20 (out_data_22_20),
		.in_data_22_21 (out_data_22_21),
		.in_data_22_22 (out_data_22_22),
		.in_data_22_23 (out_data_22_23),
		.in_data_22_24 (out_data_22_24),
		.in_data_22_25 (out_data_22_25),
		.in_data_22_26 (out_data_22_26),
		.in_data_22_27 (out_data_22_27),
		.in_data_22_28 (out_data_22_28),
		.in_data_22_29 (out_data_22_29),
		.in_data_22_30 (out_data_22_30),
		.in_data_22_31 (out_data_22_31),
		.in_data_23_0 (out_data_23_0),
		.in_data_23_1 (out_data_23_1),
		.in_data_23_2 (out_data_23_2),
		.in_data_23_3 (out_data_23_3),
		.in_data_23_4 (out_data_23_4),
		.in_data_23_5 (out_data_23_5),
		.in_data_23_6 (out_data_23_6),
		.in_data_23_7 (out_data_23_7),
		.in_data_23_8 (out_data_23_8),
		.in_data_23_9 (out_data_23_9),
		.in_data_23_10 (out_data_23_10),
		.in_data_23_11 (out_data_23_11),
		.in_data_23_12 (out_data_23_12),
		.in_data_23_13 (out_data_23_13),
		.in_data_23_14 (out_data_23_14),
		.in_data_23_15 (out_data_23_15),
		.in_data_23_16 (out_data_23_16),
		.in_data_23_17 (out_data_23_17),
		.in_data_23_18 (out_data_23_18),
		.in_data_23_19 (out_data_23_19),
		.in_data_23_20 (out_data_23_20),
		.in_data_23_21 (out_data_23_21),
		.in_data_23_22 (out_data_23_22),
		.in_data_23_23 (out_data_23_23),
		.in_data_23_24 (out_data_23_24),
		.in_data_23_25 (out_data_23_25),
		.in_data_23_26 (out_data_23_26),
		.in_data_23_27 (out_data_23_27),
		.in_data_23_28 (out_data_23_28),
		.in_data_23_29 (out_data_23_29),
		.in_data_23_30 (out_data_23_30),
		.in_data_23_31 (out_data_23_31),
		.in_data_24_0 (out_data_24_0),
		.in_data_24_1 (out_data_24_1),
		.in_data_24_2 (out_data_24_2),
		.in_data_24_3 (out_data_24_3),
		.in_data_24_4 (out_data_24_4),
		.in_data_24_5 (out_data_24_5),
		.in_data_24_6 (out_data_24_6),
		.in_data_24_7 (out_data_24_7),
		.in_data_24_8 (out_data_24_8),
		.in_data_24_9 (out_data_24_9),
		.in_data_24_10 (out_data_24_10),
		.in_data_24_11 (out_data_24_11),
		.in_data_24_12 (out_data_24_12),
		.in_data_24_13 (out_data_24_13),
		.in_data_24_14 (out_data_24_14),
		.in_data_24_15 (out_data_24_15),
		.in_data_24_16 (out_data_24_16),
		.in_data_24_17 (out_data_24_17),
		.in_data_24_18 (out_data_24_18),
		.in_data_24_19 (out_data_24_19),
		.in_data_24_20 (out_data_24_20),
		.in_data_24_21 (out_data_24_21),
		.in_data_24_22 (out_data_24_22),
		.in_data_24_23 (out_data_24_23),
		.in_data_24_24 (out_data_24_24),
		.in_data_24_25 (out_data_24_25),
		.in_data_24_26 (out_data_24_26),
		.in_data_24_27 (out_data_24_27),
		.in_data_24_28 (out_data_24_28),
		.in_data_24_29 (out_data_24_29),
		.in_data_24_30 (out_data_24_30),
		.in_data_24_31 (out_data_24_31),
		.in_data_25_0 (out_data_25_0),
		.in_data_25_1 (out_data_25_1),
		.in_data_25_2 (out_data_25_2),
		.in_data_25_3 (out_data_25_3),
		.in_data_25_4 (out_data_25_4),
		.in_data_25_5 (out_data_25_5),
		.in_data_25_6 (out_data_25_6),
		.in_data_25_7 (out_data_25_7),
		.in_data_25_8 (out_data_25_8),
		.in_data_25_9 (out_data_25_9),
		.in_data_25_10 (out_data_25_10),
		.in_data_25_11 (out_data_25_11),
		.in_data_25_12 (out_data_25_12),
		.in_data_25_13 (out_data_25_13),
		.in_data_25_14 (out_data_25_14),
		.in_data_25_15 (out_data_25_15),
		.in_data_25_16 (out_data_25_16),
		.in_data_25_17 (out_data_25_17),
		.in_data_25_18 (out_data_25_18),
		.in_data_25_19 (out_data_25_19),
		.in_data_25_20 (out_data_25_20),
		.in_data_25_21 (out_data_25_21),
		.in_data_25_22 (out_data_25_22),
		.in_data_25_23 (out_data_25_23),
		.in_data_25_24 (out_data_25_24),
		.in_data_25_25 (out_data_25_25),
		.in_data_25_26 (out_data_25_26),
		.in_data_25_27 (out_data_25_27),
		.in_data_25_28 (out_data_25_28),
		.in_data_25_29 (out_data_25_29),
		.in_data_25_30 (out_data_25_30),
		.in_data_25_31 (out_data_25_31),
		.in_data_26_0 (out_data_26_0),
		.in_data_26_1 (out_data_26_1),
		.in_data_26_2 (out_data_26_2),
		.in_data_26_3 (out_data_26_3),
		.in_data_26_4 (out_data_26_4),
		.in_data_26_5 (out_data_26_5),
		.in_data_26_6 (out_data_26_6),
		.in_data_26_7 (out_data_26_7),
		.in_data_26_8 (out_data_26_8),
		.in_data_26_9 (out_data_26_9),
		.in_data_26_10 (out_data_26_10),
		.in_data_26_11 (out_data_26_11),
		.in_data_26_12 (out_data_26_12),
		.in_data_26_13 (out_data_26_13),
		.in_data_26_14 (out_data_26_14),
		.in_data_26_15 (out_data_26_15),
		.in_data_26_16 (out_data_26_16),
		.in_data_26_17 (out_data_26_17),
		.in_data_26_18 (out_data_26_18),
		.in_data_26_19 (out_data_26_19),
		.in_data_26_20 (out_data_26_20),
		.in_data_26_21 (out_data_26_21),
		.in_data_26_22 (out_data_26_22),
		.in_data_26_23 (out_data_26_23),
		.in_data_26_24 (out_data_26_24),
		.in_data_26_25 (out_data_26_25),
		.in_data_26_26 (out_data_26_26),
		.in_data_26_27 (out_data_26_27),
		.in_data_26_28 (out_data_26_28),
		.in_data_26_29 (out_data_26_29),
		.in_data_26_30 (out_data_26_30),
		.in_data_26_31 (out_data_26_31),
		.in_data_27_0 (out_data_27_0),
		.in_data_27_1 (out_data_27_1),
		.in_data_27_2 (out_data_27_2),
		.in_data_27_3 (out_data_27_3),
		.in_data_27_4 (out_data_27_4),
		.in_data_27_5 (out_data_27_5),
		.in_data_27_6 (out_data_27_6),
		.in_data_27_7 (out_data_27_7),
		.in_data_27_8 (out_data_27_8),
		.in_data_27_9 (out_data_27_9),
		.in_data_27_10 (out_data_27_10),
		.in_data_27_11 (out_data_27_11),
		.in_data_27_12 (out_data_27_12),
		.in_data_27_13 (out_data_27_13),
		.in_data_27_14 (out_data_27_14),
		.in_data_27_15 (out_data_27_15),
		.in_data_27_16 (out_data_27_16),
		.in_data_27_17 (out_data_27_17),
		.in_data_27_18 (out_data_27_18),
		.in_data_27_19 (out_data_27_19),
		.in_data_27_20 (out_data_27_20),
		.in_data_27_21 (out_data_27_21),
		.in_data_27_22 (out_data_27_22),
		.in_data_27_23 (out_data_27_23),
		.in_data_27_24 (out_data_27_24),
		.in_data_27_25 (out_data_27_25),
		.in_data_27_26 (out_data_27_26),
		.in_data_27_27 (out_data_27_27),
		.in_data_27_28 (out_data_27_28),
		.in_data_27_29 (out_data_27_29),
		.in_data_27_30 (out_data_27_30),
		.in_data_27_31 (out_data_27_31),
		.in_data_28_0 (out_data_28_0),
		.in_data_28_1 (out_data_28_1),
		.in_data_28_2 (out_data_28_2),
		.in_data_28_3 (out_data_28_3),
		.in_data_28_4 (out_data_28_4),
		.in_data_28_5 (out_data_28_5),
		.in_data_28_6 (out_data_28_6),
		.in_data_28_7 (out_data_28_7),
		.in_data_28_8 (out_data_28_8),
		.in_data_28_9 (out_data_28_9),
		.in_data_28_10 (out_data_28_10),
		.in_data_28_11 (out_data_28_11),
		.in_data_28_12 (out_data_28_12),
		.in_data_28_13 (out_data_28_13),
		.in_data_28_14 (out_data_28_14),
		.in_data_28_15 (out_data_28_15),
		.in_data_28_16 (out_data_28_16),
		.in_data_28_17 (out_data_28_17),
		.in_data_28_18 (out_data_28_18),
		.in_data_28_19 (out_data_28_19),
		.in_data_28_20 (out_data_28_20),
		.in_data_28_21 (out_data_28_21),
		.in_data_28_22 (out_data_28_22),
		.in_data_28_23 (out_data_28_23),
		.in_data_28_24 (out_data_28_24),
		.in_data_28_25 (out_data_28_25),
		.in_data_28_26 (out_data_28_26),
		.in_data_28_27 (out_data_28_27),
		.in_data_28_28 (out_data_28_28),
		.in_data_28_29 (out_data_28_29),
		.in_data_28_30 (out_data_28_30),
		.in_data_28_31 (out_data_28_31),
		.in_data_29_0 (out_data_29_0),
		.in_data_29_1 (out_data_29_1),
		.in_data_29_2 (out_data_29_2),
		.in_data_29_3 (out_data_29_3),
		.in_data_29_4 (out_data_29_4),
		.in_data_29_5 (out_data_29_5),
		.in_data_29_6 (out_data_29_6),
		.in_data_29_7 (out_data_29_7),
		.in_data_29_8 (out_data_29_8),
		.in_data_29_9 (out_data_29_9),
		.in_data_29_10 (out_data_29_10),
		.in_data_29_11 (out_data_29_11),
		.in_data_29_12 (out_data_29_12),
		.in_data_29_13 (out_data_29_13),
		.in_data_29_14 (out_data_29_14),
		.in_data_29_15 (out_data_29_15),
		.in_data_29_16 (out_data_29_16),
		.in_data_29_17 (out_data_29_17),
		.in_data_29_18 (out_data_29_18),
		.in_data_29_19 (out_data_29_19),
		.in_data_29_20 (out_data_29_20),
		.in_data_29_21 (out_data_29_21),
		.in_data_29_22 (out_data_29_22),
		.in_data_29_23 (out_data_29_23),
		.in_data_29_24 (out_data_29_24),
		.in_data_29_25 (out_data_29_25),
		.in_data_29_26 (out_data_29_26),
		.in_data_29_27 (out_data_29_27),
		.in_data_29_28 (out_data_29_28),
		.in_data_29_29 (out_data_29_29),
		.in_data_29_30 (out_data_29_30),
		.in_data_29_31 (out_data_29_31),
		.in_data_30_0 (out_data_30_0),
		.in_data_30_1 (out_data_30_1),
		.in_data_30_2 (out_data_30_2),
		.in_data_30_3 (out_data_30_3),
		.in_data_30_4 (out_data_30_4),
		.in_data_30_5 (out_data_30_5),
		.in_data_30_6 (out_data_30_6),
		.in_data_30_7 (out_data_30_7),
		.in_data_30_8 (out_data_30_8),
		.in_data_30_9 (out_data_30_9),
		.in_data_30_10 (out_data_30_10),
		.in_data_30_11 (out_data_30_11),
		.in_data_30_12 (out_data_30_12),
		.in_data_30_13 (out_data_30_13),
		.in_data_30_14 (out_data_30_14),
		.in_data_30_15 (out_data_30_15),
		.in_data_30_16 (out_data_30_16),
		.in_data_30_17 (out_data_30_17),
		.in_data_30_18 (out_data_30_18),
		.in_data_30_19 (out_data_30_19),
		.in_data_30_20 (out_data_30_20),
		.in_data_30_21 (out_data_30_21),
		.in_data_30_22 (out_data_30_22),
		.in_data_30_23 (out_data_30_23),
		.in_data_30_24 (out_data_30_24),
		.in_data_30_25 (out_data_30_25),
		.in_data_30_26 (out_data_30_26),
		.in_data_30_27 (out_data_30_27),
		.in_data_30_28 (out_data_30_28),
		.in_data_30_29 (out_data_30_29),
		.in_data_30_30 (out_data_30_30),
		.in_data_30_31 (out_data_30_31),
		.in_data_31_0 (out_data_31_0),
		.in_data_31_1 (out_data_31_1),
		.in_data_31_2 (out_data_31_2),
		.in_data_31_3 (out_data_31_3),
		.in_data_31_4 (out_data_31_4),
		.in_data_31_5 (out_data_31_5),
		.in_data_31_6 (out_data_31_6),
		.in_data_31_7 (out_data_31_7),
		.in_data_31_8 (out_data_31_8),
		.in_data_31_9 (out_data_31_9),
		.in_data_31_10 (out_data_31_10),
		.in_data_31_11 (out_data_31_11),
		.in_data_31_12 (out_data_31_12),
		.in_data_31_13 (out_data_31_13),
		.in_data_31_14 (out_data_31_14),
		.in_data_31_15 (out_data_31_15),
		.in_data_31_16 (out_data_31_16),
		.in_data_31_17 (out_data_31_17),
		.in_data_31_18 (out_data_31_18),
		.in_data_31_19 (out_data_31_19),
		.in_data_31_20 (out_data_31_20),
		.in_data_31_21 (out_data_31_21),
		.in_data_31_22 (out_data_31_22),
		.in_data_31_23 (out_data_31_23),
		.in_data_31_24 (out_data_31_24),
		.in_data_31_25 (out_data_31_25),
		.in_data_31_26 (out_data_31_26),
		.in_data_31_27 (out_data_31_27),
		.in_data_31_28 (out_data_31_28),
		.in_data_31_29 (out_data_31_29),
		.in_data_31_30 (out_data_31_30),
		.in_data_31_31 (out_data_31_31),
		.out_data (mux_data_out)
	);

endmodule
